Särskild rapport
SMF-instrumentet i praktiken:
ett ändamålsenligt och
innovativt program som
står inför utmaningar
Innehållsförteckning
Punkt
Sammanfattning
I–XIV
Inledning
01–20
Vikten av små och medelstora företag och innovation i EU:s
ekonomi
01–03
Större fokus på små och medelstora företag och innovation i
Horisont 2020
04–06
Vad är SMF-instrumentet?
07–12
En kortfattad historik över SMF-instrumentet
13–20
Revisionens inriktning och omfattning samt
revisionsmetod
21–26
Iakttagelser
27–128
Inriktning på rätt stödmottagare
27–39
SMF-instrumentets syften och målgrupp har förändrats under dess
genomförande
28–34
Det sena införandet av konceptet icke bankmässig säkerhet
35–39
Geografisk täckning
40–58
Varierande deltagandenivåer mellan länderna – beror delvis på faktorer som
kommissionen inte kan påverka
40–49
Medvetenheten påverkades av frånvaron av en målinriktad
marknadsförings- och kommunikationsstrategi på kommissionsnivå
50–58
Urval av projekt
59–79
Begränsade utvärderingsresurser och ett distansutvärderingsförfarande som
är överbelastat på grund av ett stort antal ansökningar
61–64
Presentation inför en jury förbättrar i hög grad urvalsförfarandet samtidigt
som tiden för bidragsbeviljande hålls
65–69
Vissa it-verktyg utgör en risk för utvärderingsprocessen
70–73
Förslag som lämnas in på nytt är betungande för utvärderingsresurserna
74–79
Stödets ändamålsenlighet i SMF-instrumentets faser
80–105
Fas 1 ger användbart stöd till små och medelstora företag men det finns
redan liknande system i vissa medlemsstater
81–86
Fas 1 är alltför betungande för förvaltningen av SMF-instrumentet
87–90
Fas 2 ger ändamålsenligt stöd till små och medelstora företag
91–94
Företagsaccelerationstjänsterna i fas 3 har potential, men de lanserades
sent
95–103
SMF-instrumentets ändamålsenlighet har inte bedömts, och dess framtida
roll i Horisont Europa har ännu inte fastställts
104–105
Locka till sig investeringar efter finansieringen genom SMFinstrumentet
106–128
Kommissionen har bara begränsad kunskap om stödmottagarnas
övergripande finansieringsbehov och har inte skapat länkar till EU:s
finansieringsinstrument
107–116
Stödmottagarna lockar till sig ytterligare investeringar, men nivåerna
varierar i EU
117–128
Slutsatser och rekommendationer
129–139
Inriktning på rätt stödmottagare
Geografisk täckning
Urval av projekt
133–135
Stödets ändamålsenlighet i SMF-instrumentets faser
136–138
Locka till sig investeringar efter finansieringen genom SMF-instrumentet
Bilagor
Bilaga I – Metod
Bilaga II – Statistik
Bilaga III – Europeiska innovationsrådet inom ramen för
Horisont Europa – från idé till förslag
Akronymer och förkortningar
Ordlista
Kommissionens svar
Granskningsteam
Tidslinje
Sammanfattning
I Instrumentet för små och medelstora företag inrättades genom ramprogrammet för
forskning, Horisont 2020, för att stödja innovation i små eller medelstora företag
(SMF). Syftet är att utveckla och utnyttja potentialen hos små och medelstora företag
genom att avhjälpa bristen på finansiering för nystartade projekt med hög risk och öka
den privata kommersialiseringen av forskningsresultat. Instrumentet riktar sig till
innovativa små och medelstora företag i EU och 16 associerade länder som visar en
stark strävan att utvecklas, växa och internationaliseras genom alla olika typer av
innovation.
II Med en sammanlagd budget på 3 miljarder euro för perioden 2014–2020 beviljar
instrumentet bidrag till företag med stor potential, för att stödja dem antingen i
utarbetandet av en genomförbarhetsstudie (upp till 50 000 euro i fas 1) eller i
samband med deras forskning och utveckling och marknadstester (2,5 miljoner euro i
fas 2). Stöd kan också ges i form av coachning, mentorskap eller andra tjänster för
företagsacceleration (fas 3).
III I denna revision utvärderade vi huruvida SMF-instrumentet stöder innovation i
små och medelstora företag. Vi undersökte om instrumentet har riktat in sig på rätt
typ av små och medelstora företag, om det uppnådde en bred geografisk täckning, om
urvalsförfarandet och stödet från kommissionen var ändamålsenligt och om
kommissionen övervakade och följde upp instrumentet på rätt sätt för att
åstadkomma förbättringar. Vi förväntar oss att våra iakttagelser och de
rekommendationer som vi gör används som underlag i diskussionen om hur SMFinstrumentets efterträdare ska inrättas och förvaltas efter 2020 och framåt.
IV Vi konstaterade att SMF-instrumentet ger ett ändamålsenligt stöd till små och
medelstora företag när de utvecklar sina innovationsprojekt och att det EU-varumärke
som följer av EU-stödet hjälper företagen att locka till sig ytterligare investeringar.
V Instrumentets breda syften och mål har dock, tillsammans med de ändringar som
gjorts under genomförandet, skapat ovisshet bland intressenterna. Vi konstaterade att
det finns en risk för att instrumentet finansierar vissa små och medelstora företag som
skulle ha kunnat få finansiering på marknaden.
VI Deltagandet i SMF-instrumentet varierar stort mellan medlemsstaterna. Detta
beror till viss del på externa faktorer men också på de varierande nivåer av stöd som
tillhandahålls av nationella kontaktpunkter och på begränsningar i fråga om
kommissionens marknadsförings- och kommunikationsverksamhet.
VII Vi konstaterade att utvärderings- och urvalsförfarandena har förbättrats under
instrumentets livstid. Den muntliga presentationen av projektförslag inför en panel av
jurymedlemmar bidrar på ett särskilt värdefullt sätt till urvalet av de bästa förslagen.
Det saknas dock ömsesidig återkoppling mellan utvärderingsstegen. Dessutom är vissa
it-verktyg inte ändamålsenliga, vilket påverkar en redan pressad process negativt.
VIII Att förslag som tidigare inte valts ut lämnas in på nytt är en stor och allt större
belastning för förvaltnings- och utvärderingsresurserna, som inte tillför något
mervärde. Detta ökar inte bara de administrativa kostnaderna utan sänker också
framgångsgraden, det vill säga andelen ansökningar som beviljas stöd, och avskräcker
på så sätt företag från att delta.
IX Instrumentets fas 1 tillhandahåller ändamålsenligt stöd tack vare sin enkla och
snabba urvalsprocess, EU:s varumärke och tillgången till företagsaccelerationstjänster.
Denna fas innebär dock oproportionerligt höga administrativa kostnader för
kommissionens förvaltning, och instrumentets relevans minskar i länder där det redan
finns liknande program.
X Fas 2 av instrumentet, som ger en högre nivå av stöd med målet att lansera
innovationen på marknaden, har samma positiva utfall som fas 1 och hjälper också
små och medelstora företag att dra till sig ytterligare investeringar.
XI Vi konstaterade trots detta att majoriteten av stödmottagarna fortfarande
behöver ytterligare finansiering för att stödja sitt innovationsarbete och lansera sina
projekt på marknaden. Kommissionen har inte gjort mycket för att skapa kopplingar
mellan de små och medelstora företagens finansieringsbehov och EU-stödda
finansieringsinstrument och har begränsad kunskap om stödmottagarnas behov av
finansiering.
XII Tjänsterna för coachning och företagsacceleration har potential att stärka
instrumentets effekter, men eftersom de lanserades sent var det bara ett fåtal små och
medelstora företag som använde sig av dem. De har inte heller varit tillräckligt
anpassade efter stödmottagarnas behov.
XIII Övervakningen av de investeringar som anskaffats och företagsutvecklingen är
kostnadseffektiv men bedömer inte instrumentets verkliga effekter. Även om
stödmottagarna har lyckats anskaffa investeringar utöver de bidrag som erhållits, råder
det fortfarande obalans mellan de länder som deltar: små och medelstora företag i
nordvästra Europa anskaffar mer privat finansiering än sådana företag i södra och
östra Europa.
XIV I rapporten rekommenderar vi att kommissionen gör följande:
—
Förbättrar instrumentets marknadsförings- och kommunikationsstrategi.
—
Förbättrar sitt stöd till de nationella kontaktpunkterna för små och medelstora
företag liksom till Enterprise Europe Network (EEN) och anpassar instrumentets
urvalsförfarande för att dra bättre nytta av resurserna och finansiera de bästa
förslagen.
—
Begränsar antalet gånger ett förslag får lämnas in på nytt och offentliggör
framgångsgraden per projektförslag.
—
Föreslår för medlemsstaterna att kommissionen ska förvalta system som liknar
fas 1.
—
Behåller ett system som liknar fas 2 under nästa programperiod och utgår från de
befintliga resultaten.
—
Förbättrar företagsaccelerationstjänsterna genom att tilldela lämpliga resurser.
—
Identifierar och främjar synergier mellan SMF-instrumentet och EU-stödda
finansieringsinstrument.
Inledning
Vikten av små och medelstora företag och innovation i EU:s
ekonomi
Enligt Europeiska kommissionens årsrapport om små och medelstora företag
2017/2018 utgör dessa företag 99 % av alla företag som är verksamma i EU:s ickefinansiella affärssektor, och står för 66 % av den totala sysselsättningen och 57 % av
mervärdet inom EU:s icke-finansiella affärssektor.
Både Europaparlamentet och rådet har betonat vikten av att stödja innovation (i
synnerhet banbrytande innovation) och tillväxt hos uppstartsföretag och små och
medelstora företag. De har noterat att stöd till innovativa små och medelstora företag
och uppstartsföretag är avgörande för att maximera Europas potential för tillväxt och
socioekonomisk omvandling 1. Akademiska studier 2,3 har visat på kopplingen mellan
företagande, verksamheten i små och medelstora företag, ekonomisk tillväxt och
skapande av sysselsättning.
Europa 2020-strategin4 understryker betydelsen av innovation när det gäller att
stärka EU:s tillväxt och sysselsättning. ”Innovationsunionen” är en av unionens sju
flaggskeppsinitiativ, som syftar till att skapa en innovationsvänlig miljö för att det ska
bli lättare för innovativa idéer att omvandlas till produkter och tjänster som skapar
tillväxt och arbetstillfällen 5.
Konsekvensbedömning av EU:s nionde ramprogram för forskning och innovation (en ny
horisont för Europa).
The vital 6 per cent. How high-growth innovative businesses generate prosperity and jobs
– Nesta (National Endowment for Science, Technology and the Arts).
Henrekson, M. & Johansson, D. 2010. ”Gazelles as job creators: a survey and interpretation
of the evidence”, Small Business Economics, 35, 227–244, s. 240.
Kommissionens meddelande Europa 2020 – En strategi för smart och hållbar tillväxt för alla
(KOM(2010) 2020 slutlig).
https://ec.europa.eu/info/research-and-innovation/strategy/goals-research-andinnovation-policy/innovation-uni
Större fokus på små och medelstora företag och innovation i
Horisont 2020
Horisont 2020 är EU:s åttonde ramprogram för forskning. Med en budget på
76,4 miljarder euro för perioden 2014–2020 är det världens största offentliga
forsknings- och innovationsprogram 6.
Horisont 2020 har fokuserat mer på innovation än något av de tidigare
programmen genom att tillhandahålla mer finansiering för testning,
prototypframställning, affärsdriven FoU och främjande av innovativt entreprenörskap.
Horisont 2020 har också fastställt ett mer ambitiöst mål för de medel som ska tilldelas
små och medelstora företag än något annat tidigare ramprogram: Små och medelstora
företag bör erhålla minst 20 % av den totala sammanlagda budgeten på 9 miljarder
euro inom ramen för pelarna ”Ledarskap inom möjliggörande teknik och
industriteknik” och ”Samhällsutmaningar”.
En budget på 3 miljarder euro har öronmärkts för SMF-instrumentet (SMF-I),
vilket motsvarar 33 % av SMF-målet för hela Horisont 2020 7.
Vad är SMF-instrumentet?
Instrumentet för små och medelstora företag (SMF-I) inrättades genom
ramprogrammet för forskning, Horisont 2020, för att stödja innovation i små eller
medelstora företag. Det beviljar bidrag till företag med stor potential att stödja dem i
utarbetandet av en genomförbarhetsstudie (fas 1) och i samband med deras forskning
och utveckling (FoU) och marknadstester (fas 2). Stöd kan också ges i form av
coachning, mentorskap eller andra tjänster för företagsacceleration (fas 3). SMF-I är
tillgängligt för små och medelstora företag i medlemsstaterna och i länder som har
tecknat ett associeringsavtal (associerade länder)8, och har som mål att hjälpa företag
att expandera och internationaliseras.
Förordning (EU) nr 1291/2013 om inrättande av Horisont 2020.
Förordning (EU) nr 1291/2013.
http://ec.europa.eu/research/bitlys/h2020_associated_countries.html
SMF-I är ett nytt instrument på så sätt att det låter små och medelstora företag
delta som enskilda stödmottagare utan att nödvändigtvis ingå i ett konsortium, vilket
ramprogrammen för forskning vanligtvis kräver. Det riktar sig till projekt som redan har
uppnått åtminstone nivå 6 vad gäller teknisk mognadsgrad.
Syftet med SMF-I är att utveckla och utnyttja potentialen hos små och medelstora
företag, genom att avhjälpa bristen på finansiering för nystartade forsknings- och
innovationsprojekt med hög risk och öka den privata kommersialiseringen av
forskningsresultat. Instrumentet riktar sig till små och medelstora företag som visar en
stark strävan att utvecklas, växa och internationaliseras, och ska erbjudas för alla typer
av innovation där varje verksamhet har ett tydligt europeiskt mervärde.
Det är kommissionens generaldirektorat för forskning och innovation som
ansvarar för den politiska utvecklingen av SMF-I, men instrumentet genomförs av
Genomförandeorganet för små och medelstora företag (Easme).
Instrumentet är uppdelat i tre faser (se figur 1):
—
Fas 1 (utredning av den tekniska och kommersiella genomförbarheten hos
en affärsidé): Stöd till att undersöka om en ny idé är vetenskapligt och
tekniskt genomförbar och om den har kommersiell potential. Bidrag på
euro beviljas med en medfinansieringsgrad från EU på 70 %.
—
Fas 2 (utveckling och demonstration): Utveckling av innovation i
demonstrationssyfte, prestationskontroll, provning, utveckling av
pilotverksamhet, validering inför marknadsintroduktion och annan
verksamhet som syftar till att göra innovationer investeringsberedda och
tillräckligt mogna för marknadsetablering. Bidrag på upp till 2,5 miljoner euro
kan beviljas med en medfinansieringsgrad på 70 %.
—
Fas 3 (ytterligare EU-stöd för att ta sig in på marknaden): Tillhandahållande
av stöd, utbildning och coachning, liksom underlättad tillgång till
riskfinansiering. Denna fas består av en kombination av de olika tjänster som
erbjuds stödmottagarna i faserna 1 och 2. Inga ytterligare bidrag beviljas i
denna fas.
Trots att de olika faserna är numrerade är SMF-I inte ett instrument som
genomförs i en följd: Man måste alltså inte ha genomgått fas 1 för att kunna delta i
fas 2. De tjänster som erbjuds i fas 3 kan tillhandahållas när som helst under
genomförandet av innovationsprojektet, till och med när det har slutförts.
Figur 1 – SMF-I: Struktur och budgetfördelning
SMF-I, BUDGETFÖRDELNING
Från idé till koncept
Engångsbelopp om 50 000 euro
Sex månaders genomförande
Utfall: genomförbarhetsstudie
~88 %
 Från koncept till
marknadsmognad
 Bidrag från 0,5 till 2,5 milj. euro
 Upp till 70 % av de stödberättigande
kostnaderna
 24 månaders genomförande
 Utfall: innovativ produkt, process
eller tjänst som är färdig för
marknaden
2014–maj 2019
projekt
milj. euro
projekt
FAS 2
Fas 2
2014–maj 2019
~7 %
Fas 1




~2 %
milj. euro
FAS 1
Fas 3
FAS 3
 Företagsacceleration: mässor,
förmedlingsevenemang, matchning med investerare etc.
 Coachning: tillhandahålls av EEN-utvalda coacher
~3 % – övriga utgifter
Källa: Revisionsrätten.
En kortfattad historik över SMF-instrumentet
SMF-instrumentet lanserades 2014 och utformades med utgångspunkt i USA:s
SBIR 9-program. Genom ”trattmodellen” skulle man göra ett stort antal mindre
investeringar i genomförbarhetsstudier för lovande innovationsprojekt (fas 1), där de
bästa skulle gå vidare till fas 2 och få mer finansiering. Skyldigheten att genomgå fas 1
före fas 2 ströks dock under utarbetandet och gjorde det möjligt för sökande att
ansöka direkt till vilkendera.
I likhet med andra delar av Horisont 2020 genomförs SMF-instrumentet genom
arbetsprogram, som löper över två eller tre år. Med varje arbetsprogram kan
instrumentets egenskaper ändras utifrån de politiska ambitionerna.
Arbetsprogrammen under 2014–2015 och 2016–2017 delade in budgeten för
SMF-I i olika tematiska ämnen, till exempel bioteknik, hälso- och sjukvård och säkerhet.
Små och medelstora företag skulle ansöka till det ämne som passade deras projekt
bäst.
https://www.sbir.gov/about/about-sbir
Arbetsprogrammet för 2018–2020 innehöll initiativet ”pilotprojektet för ett
europeiskt innovationsråd”, som grupperade SMF-I tillsammans med vissa andra
program – framtida framväxande teknik (FET Open), snabbspåret till innovation (FTI)
och Horisont 2020-priserna. Följande huvudsakliga ändringar som infördes under
pilotprojektet påverkade SMF-I:
o
En bottom-up-strategi med öppen ansökningsomgång utan att företagen behövde
ansöka till ett tematiskt ämne.
o
Kravet på att företagen skulle hålla en presentation för att väljas ut i fas 2:
personliga intervjuer med en panel av erfarna innovatörer.
o
Utökade möjligheter till mentorskap och coachning för alla stödmottagare under
fas 3.
I juni 2018 lade kommissionen fram ett förslag till en förordning om inrättande av
Horisont Europa för perioden efter 2020 10. I förslaget planeras ett
europeiskt innovationsråd (EIC) som den tredje pelaren i ett ramprogram med en
budget på 10,5 miljarder euro som skulle samla allt EU-stöd till banbrytande
innovation som skapar nya marknader på ett ställe och omfatta två instrument:
Pathfinder för avancerad forskning och Accelerator. Därmed skulle den tidigare fas 1
slutgiltigt läggas ner, medan åtgärder som liknar de under de tidigare fas 2 och fas 3
skulle inkluderas i Accelerator 11.
COM(2018) 435, Förslag till förordning om inrättande av Horisont Europa, juni 2018.
I april 2019 nådde kommissionen, Europaparlamentet och rådet en preliminär
överenskommelse om Horisont Europa.
I mars 2019 ändrade kommissionen arbetsprogrammet och lanserade det
utökade pilotprojektet för ett europeiskt innovationsråd, som ska löpa mellan juni
och slutet av 2020. Detta utökade projekt utgör en övergång mot det föreslagna
Europeiska innovationsrådet inom ramen för Horisont Europa (efter 2020). Det ska
skapa närmare kopplingar mellan de ingående delarna och innebär betydande
ändringar av SMF-I. Fas 1 lades ner och följande instrument lanserades:
o
Pathfinder”, som ersätter FET-Open och FET-Proactive.
o
Accelerator”, som ersätter fas 2:
—
Utveckling och uppskalning av högriskinnovation i små och medelstora
företag.
—
Införande av konceptet icke bankmässig säkerhet 12.
—
Bidrag på upp till 2,5 miljoner euro.
—
Möjlighet till kapitaltillskott på upp till 15 miljoner euro (blandad
finansiering).
Europeiska innovationsrådets pilotprojekt var en utveckling av SMF-I, som till
största delen var i linje med instrumentets ursprungliga utformning. Det utökade
pilotprojektet införde även ändringar för att underlätta en övergång till det föreslagna
europeiska innovationsrådet inom ramen för Horisont Europa. SMF-I är den största
delen av både pilotprojektet och det utökade pilotprojektet, och står för omkring två
tredjedelar av deras respektive budgetar.
Förslaget om inrättande av ett europeiskt innovationsråd genom
Horisont Europa, som för närvarande befinner sig i lagstiftningsfasen, behåller vissa av
instrumentets delar, till exempel fortsatt fokus på små och medelstora företag och
stöd som uteslutande tar formen av bidrag. Vissa andra aspekter som övervägs måste
dock fortfarande utvecklas eller testas 13.
Konceptet icke bankmässig säkerhet definieras i vanliga frågor till Europeiska
innovationsrådet som oförmåga att attrahera tillräcklig finansiering.
Till exempel tillhandahållande av ekonomiskt stöd till projekt genom finansiering med eget
kapital, och att man till viss del kan godta urvalsförfaranden som utförs i andra
ansökningsomgångar eller program.
Revisionens inriktning och omfattning
samt revisionsmetod
Denna särskilda rapport är den senaste i en serie publikationer från
Europeiska revisionsrätten som granskar ekonomiskt stöd till innovativa små och
medelstora företag14. Både Europaparlamentet och rådet har betonat vikten av att
stödja innovativa små och medelstora företag och uppstartsföretag för att maximera
Europas tillväxtpotential. Vi förväntar oss att de iakttagelser som följer av vår revision
och de rekommendationer som vi gör används som underlag för diskussionen om den
fleråriga budgetramen och om hur SMF-instrumentets efterträdare ska inrättas och
förvaltas efter 2020 och framåt.
I denna revision granskade vi huruvida SMF-instrumentet var ändamålsenligt när
det gäller att stödja innovation i små och medelstora företag.
I revisionen tittade vi på huruvida
o
instrumentet riktade sig till ”rätt små och medelstora företag” (dvs. sådana med
stor innovationspotential),
o
instrumentet uppnådde geografisk täckning och letade efter spetskompetens,
o
kommissionens urvalsförfarande hade utformats för att finansiera de bästa
projekten,
o
kommissionen gav stödmottagarna ändamålsenligt stöd,
o
kommissionen övervakade och följde upp instrumentet på lämpligt sätt för att
åstadkomma förbättringar.
Vår revision var därför inriktad på instrumentets utformning, förvaltning och
output, liksom dess utveckling mot ett europeiskt innovationsråd, inklusive
pilotprojektet för detta. I vår revision inkluderade vi de bidrag som beviljats mellan
januari 2014 och maj 2019.
De särskilda rapporterna om garantier (SR 20/2017 om garantiinstrumentet för små och
medelstora företag) och om riskkapital (SR 17/2019).
Revisionen kombinerade bevis från en mängd olika källor:
o
En skrivbordsgranskning av dokument.
o
En granskning av analytiska data.
o
Enkätundersökningar bland stödmottagare, icke utvalda sökande som erhållit en
spetskompetensstämpel, distansutvärderare och nationella
innovationsmyndigheter.
o
Informationsbesök i Bulgarien, Danmark, Frankrike, Rumänien, Slovenien, Spanien
och Förenade kungariket.
o
Intervjuer med kommissionens generaldirektorat, Easme,
Europeiska investeringsbanken (EIB), Europeiska investeringsfonden (EIF) och
andra berörda intressenter.
Se bilaga I för närmare uppgifter om vår revisionsmetod och våra beviskällor.
Iakttagelser
Inriktning på rätt stödmottagare
Enligt Horisont 2020-förordningen15 riktar sig SMF-I till innovativa små och
medelstora företag med en stark strävan att utvecklas, växa och internationaliseras.
SMF-instrumentets syften och målgrupp har förändrats under dess
genomförande
Instrumentets intressenter påpekade i intervjuer och svar på våra enkäter att
SMF-I skulle ha vunnit på om dess mål och syften hade definierats på ett tydligare sätt
när instrumentet togs fram.
Denna tvetydighet, i synnerhet när det gäller vilken typ av företag som
instrumentet riktade sig till, belystes också i rapporten från den rådgivande gruppen av
SMF-experter (EAG) 2014 16. Enligt EAG skulle ytterligare resurser och en mer
djupgående analys av den avsedda målgruppen ha gjort att kommissionen med större
säkerhet kunnat locka till sig rätt typ av sökande.
De efterföljande arbetsprogrammens syften förändrades flera gånger under
genomförandet. De två första arbetsprogrammen (2014–2015 och 2016–2017)
fokuserade på all slags innovation som främjande företagstillväxt och var ny för
marknaden. Arbetsprogrammet för pilotprojektet för ett europeiskt innovationsråd
(2018–2020) och det utökade pilotprojektet för ett europeiskt innovationsråd (2019–
2020) ändrade fokus mot innovation som är ”marknadsskapande”. Som en jämförelse
har SBIR-programmet inte förändrats särskilt mycket sedan det förlängdes 2011 17.
De många ändringar som gjorts under den korta tid som SMF-I har varit igång har
skapat förvirring för huvudaktörerna, bland dessa de nationella kontaktpunkterna,
Enterprise Europe Network (EEN) och de sökande, när det gäller vad som ska
finansieras.
Förordning (EU) nr 1291/2013 om inrättande av Horisont 2020.
års rapport från EAG om innovation i små och medelstora företag.
https://sbir.nih.gov/reauthorization#eligibilityDiv
Under genomförandet av SMF-I ändrades den typ av företag som instrumentet
riktade sig till, från mogna företag som hade deltagit i tidigare ramprogram till
innovativa och, i synnerhet, unga företag utan tidigare erfarenhet från ramprogram.
Införandet under 2018 av bottom-up-strategin och presentationsdelen i pilotprojektet
skyndade på en ”föryngring” bland de små och medelstora företagen (se figur 2).
Figur 2 – Ålder på små och medelstora företag som finansierats i fas 2
per ansökningsår
%
%
%
%
%
≥ 20
%
10–19
5–9
%
<5
%
%
%
0%
Källa: Revisionsrätten, på grundval av uppgifter från kommissionen.
Den nuvarande åldersprofilen bland stödmottagarna matchar den för de företag
som identifierades i Nesta-studien 18 om företags tillväxtfaktorer och skillnader i
skapandet av arbetstillfällen. Detta visar att den nuvarande uppsättningen
stödmottagare har bättre möjlighet att generera tillväxt och skapa arbetstillfällen.
Bottom-up-strategin har löst problemet med den tidigare strukturen där
företagen kunde välja att söka stöd inom ett visst ”ämne” baserat på skillnader i
framgångsgrad. Den har också förenklat ansökningsomgångarnas administrativa
förfaranden. En alternativ strategi kan vara lämplig i de fall det finns ett behov att
öronmärka specifika områden som anses prioriterade för EU.
Arbetsdokument från Nesta nr 11/02, A look at business growth and contraction in Europe.
Det sena införandet av konceptet icke bankmässig säkerhet
SMF-I syftar till att ”avhjälpa bristen på finansiering av inledande forskning och
innovation med hög risk” 19. De efterföljande arbetsprogrammen har dock inte
specificerat hur man ska nå små och medelstora företag som har svårt att erhålla
finansiering från andra källor, och konceptet icke bankmässig säkerhet infördes först
genom det utökade pilotprojektet för ett europeiskt innovationsråd under 2019.
Enligt flera intressenter som intervjuades finns det en risk för att SMF-I tränger ut
privata investeringar. Denna slutsats kunde dras från resultatet av den enkät som vi
skickade till stödmottagare. I fas 2 trodde 36 % av de som svarade att deras projekt
skulle ha kunnat få finansiering från den privata sektorn, och 17 % svarade att de hade
kunnat använda företagets egna medel för att finansiera innovationen.
Jurymedlemmarna bekräftade också denna risk i intervjuer (se figur 3).
Figur 3 – Fas 2-företags alternativa källor till privat finansiering
0%
%
%
%
%
%
Privat sektor
Egna medel
Ja
Nej
Vet ej
Källa: Revisionsrättens enkät till stödmottagare.
Intressenterna framhöll dock den efterföljande förstärkningseffekt som uppstod
på grund av EU-bidraget och som hjälper stödmottagarna att senare attrahera de
ytterligare medel som behövs för att vidareutveckla deras innovationsprojekt och
expandera.
Förordning (EU) nr 1291/2013 om inrättande av Horisont 2020.
Ett projekts bankmässiga säkerhet är ett komplext koncept som påverkas av flera
olika variabler, däribland den finansieringsvolym som behövs, tidpunkten och priset.
Med tanke på konceptets komplexa karaktär ansåg de flesta som intervjuades att man
behöver definiera vad som avses med bankmässig säkerhet och hur detta ska mätas.
Före 2019 tog man inte hänsyn till projektens bankmässiga säkerhet i
urvalsförfarandena till SMF-I. Instrumentet beviljade bidrag till vissa små och
medelstora företag som skulle ha kunnat finansieras av marknaden. Införandet av
konceptet icke bankmässig säkerhet kräver tydliga regler för hur detta kan bevisas, i
synnerhet eftersom EU-varumärket som erhålls genom SMF-I och bidraget i sig lockar
till sig ytterligare finansiella resurser till stöd för stödmottagarnas innovationsprojekt.
Geografisk täckning
Varierande deltagandenivåer mellan länderna – beror delvis på faktorer
som kommissionen inte kan påverka
Spetskompetens är i högsta grad avgörande för deltagandet i SMF-I och
projektens framgång. Med tanke på de olikartade innovationsnivåerna bland
medlemsstaterna kan man därför förvänta sig att medlen fördelas ojämnt. Samtidigt
strävar dock EU, genom Horisont 2020, efter att se till att fördelarna med en
innovationsdriven ekonomi maximeras och sprids vida omkring 20.
Skäl 14 i rådets beslut 2013/743/EU.
Graferna och kartorna nedan (figur 4, bild 1 och bild 2) illustrerar statistiken på
landsnivå i fråga om antalet inlämnande förslag och den finansiering som erhållits i
förhållande till antalet små och medelstora företag, BNP och befolkning. Bilaga II visar
fördelningen av SMF-I-finansiering per medlemsstat i absoluta och relativa termer,
antalet projekt som valts ut, antalet förslag och framgångsgraden per medlemsstat.
Traditionellt sett har genomförandeanalyserna av Horisont 2020 framhållit två
olika medlemsstatsgrupper: EU-15 och EU-13 21. När det gäller SMF-instrumentet kan
denna åtskillnad inte förklara skillnaderna i den finansiering som erhållits (se den
första kolumnen i figur 4).
Figur 4 – Fördelning av SMF-I-finansiering i förhållande till antalet små
och medelstora företag, BNP och befolkning
Finansiering från SMF-I (i euro)/antal SMF
Finansiering från SMF-I (i euro)/BNP (i miljoner euro)
Danmark
Finland
Irland
Österrike
Slovenien
Österrike
Spanien
Förenade kungariket
Malta
Malta
Slovenien
Österrike
Spanien
Nederländerna
Förenade
kungariket
Malta
Tyskland
Estland
Sverige
Nederländerna
Förenade
kungariket
Tyskland
Spanien
Nederländerna
Irland
Sverige
Finland
Estland
Sverige
Slovenien
Danmark
Finland
Irland
Estland
Finansiering från SMF-I (i euro)/befolkning
Danmark
Tyskland
Frankrike
Frankrike
Frankrike
Belgien
Belgien
Belgien
Ungern
Italien
Ungern
Italien
Portugal
Litauen
Italien
Portugal
Ungern
Polen
Polen
Grekland
Grekland
Lettland
Lettland
Kroatien
Luxemburg
Cypern
Cypern
Luxemburg
Cypern
Tjeckien
Tjeckien
Bulgarien
Bulgarien
Slovakien
Rumänien
-
Slovakien
-
Kroatien
Tjeckien
Slovakien
Lettland
Bulgarien
Rumänien
Grekland
Polen
Kroatien
Litauen
Luxemburg
Portugal
Litauen
Rumänien
-
Källa: Revisionsrätten, på grundval av uppgifter från kommissionen.
Med EU-13 avses Bulgarien, Cypern, Estland, Kroatien, Lettland, Litauen, Malta, Polen,
Rumänien, Slovakien, Slovenien, Tjeckien och Ungern, medan EU-15 är de resterande 15
medlemsstaterna i Europeiska unionen.
Bild 1 – Antal inlämnade projektförslag per tusen små och medelstora
företag
Källa: Revisionsrätten.
Bild 2 – SMF-I-finansiering per SMF (i euro/SMF)
Källa: Revisionsrätten.
Deltagandenivån för SMF-I och projektens framgångsgrad påverkas av flera
faktorer:
Innovationsekosystemen och antalet små och medelstora företag i landet.
Om det finns en nationell strategi för SMF-I eller inte.
Det arbete som gjorts för att marknadsföra SMF-I.
Stödet från nationella kontaktpunkter och EEN.
Även om kommissionen inte kan påverka vissa av dessa faktorer kan den påverka
andra – såsom marknadsföringen och främjandet av instrumentet eller det stöd som
ges av de nationella kontaktpunkterna.
Skillnaderna i framgångsgrad mellan länderna kan delvis förklaras med hjälp av
den befintliga variationen i innovationsnivå. Figur 5 visar ett starkt samband mellan
framgångsgraderna i SMF-I och den europeiska resultattavlan för innovations
sammanfattande innovationsindex22.
Figur 5 – Samband mellan framgångsgraden avseende SMF-I och den
europeiska resultattavlan för innovation 2019
Europeiska resultattavlan för innovation
0,8
LU
0,6
0,5
EL
CZ
0,4
MT
CY
HU
PL
LV
0,3
BG
0,2
HR
DK
NL
UK
DE
BE
EE
SK
0,1
SE
FI
0,7
AT
IE
FR
PT
SL
it
5%
6%
7%
8%
Framgångsgrad per land
LT
ES
RO
1%
2%
3%
4%
9%
%
%
%
%
Källa: Revisionsrätten, på grundval av uppgifter från kommissionen.
https://ec.europa.eu/growth/industry/innovation/facts-figures/scoreboards_sv
Ett gemensamt drag hos deltagarländer med ett högt deltagande och höga
framgångsgrader med avseende på instrumentet är att det finns en aktiv nationell
innovationsmyndighet, som fungerar som en mellanhand för innovativa små och
medelstora företag. I de tre medlemsstater som hade lägst deltagande (jämfört med
antalet små och medelstora företag i landet) och de lägsta framgångsgraderna finns
det däremot ingen sådan myndighet.
I vår enkät till nationella innovationsmyndigheter frågade vi om de hade
nationella program där man gav stöd till små och medelstora företag som ville ansöka
till SMF-I. Knappt hälften av myndigheterna bekräftade att de hade nationella program
för stöd till små och medelstora företag som ansöker till fas 2, och 35 % rapporterade
detta för fas 1 (se figur 6). Intervjuobjekten noterade att sedan SMF-I skapades hade
vissa nationella myndigheter dragit ner på liknande program och i stället förberett
företagen för SMF-I.
Figur 6 – Finns det nationella program för stöd till små och medelstora
företag när de ansöker till fas 1 och/eller fas 2 i ert land?
Fas 1
Fas 2
0%
%
%
Ja
%
%
Nej
Källa: Revisionsrättens enkät till nationella innovationsmyndigheter.
Spanien är ett bra exempel på en medlemsstat med en nationell strategi som ger
stöd till innovativa företag som skulle kunna ansöka till SMF-I. De spanska
myndigheterna har inrättat ett system för att marknadsföra SMF-I, och letar aktivt
efter mycket innovativa företag och ger dem stöd när de ansöker till instrumentet.
Spanien är SMF-I:s största stödmottagare: landet får 20 % av den sammanlagda
budgeten och har det högsta antalet ansökande små och medelstora företag. Trots att
Spanien är en blygsam innovatör enligt den europeiska resultattavlan för innovation
har landet en av de högsta framgångsgraderna. Irland och Danmark marknadsför också
aktivt instrumentet och förbereder sina små och medelstora företag för att delta.
I de medlemsstater som besöktes och som hade ett lågt deltagande i SMF-I (vad
gäller tilldelade medel och framgångsgrad) var medvetenheten om SMF-I begränsad.
Specifikt stöd eller marknadsföring på nationell nivå, eller vägledning för företag om
instrumentet, var ovanligt. De låga framgångsgraderna har i sin tur avskräckt andra
företag från att ansöka till SMF-I. Dessutom har förekomsten av alternativa nationella
program, med högre framgångsgrader, minskat attraktionskraften för SMF-I för företag
och fristående experter, exempelvis konsulter.
Medvetenheten påverkades av frånvaron av en målinriktad
marknadsförings- och kommunikationsstrategi på kommissionsnivå
SMF-I utgör en ny form av stöd i ramprogrammen, som främst riktar sig till
enskilda små och medelstora företag med mycket innovativa projekt, med en
marknadsdriven strategi.
Traditionella Horisont 2020-sökande (universitet, stora bolag och
forskningscentrum) känner till de finansieringsmöjligheter som erbjuds genom
Horisont 2020. Dessa organisationer har erfarenhet av både Horisont 2020 och tidigare
ramprogram, och i många fall har de särskild personal som sköter ansökningar och
projekt. Den typ av företag som SMF-I riktar sig till har i regel inte deltagit i några
tidigare ramprogram och har kanske inte ens inkluderat offentliga medel i sin
finansstrategi.
Vi undersökte huruvida SMF-I marknadsfördes, genomfördes och övervakades för
att ge små och medelstora företag enkel tillgång till instrumentet, i enlighet med
rådets beslut 2013/743/EU. Vi tittade också på i vilken utsträckning
marknadsföringstekniker användes för att göra rätt företag medvetna om att denna
finansieringsmöjlighet finns, och i vilken utsträckning lämpliga kommunikationskanaler
måste identifieras och användas för att nå dem.
Kommissionen och Easme hade en begränsad budget för sin
kommunikationsverksamhet och för att anordna olika evenemang som samlade
potentiella stödmottagare inom SMF-I, främst informationsdagar för Horisont 2020.
Rapporter från EAG belyste att det saknades en marknadsföringsstrategi för SMF-I, och
att man behövde identifiera rätt ”klienter” och anpassa kommunikationskanalerna och
kommunikationsverktygen efter dessa. I utvärderingen av SMF-I 23 sågs detta som en
möjlig förklaring till de olika genomslagsgraderna i EU-28, och den pekade på behovet
av att granska kommunikations- och marknadsföringsstrategin på nytt.
Även om ansträngningar gjordes för att nå potentiella stödmottagare hade
kommissionen inte någon strukturerad marknadsförings- och kommunikationsstrategi.
Kommissionen använde inte en tillräckligt målinriktad metod för att öka
medvetenheten bland innovativa små och medelstora företag om de möjligheter som
SMF-I erbjuder.
Kommissionen förlitar sig i hög grad på den marknadsföring som sköts av de
nationella kontaktpunkterna och EEN för att uppnå ett enhetligt genomförande av
SMF-I. Den anser att kontaktpunkterna är ”den huvudsakliga strukturen för att förse
potentiella deltagare med praktisk information och hjälp”. Eftersom små och
medelstora företag är mindre bekanta med Horisont 2020 än andra deltagare i
ramprogrammet (se punkt 51) är de nationella kontaktpunkternas roll särskilt viktig för
små och medelstora företag. De nationella kontaktpunkterna utses och får betalt av de
nationella myndigheterna. De ansvarar för att säkerställa att alla potentiella sökande
blir medvetna om det nya programmet och att det blir lättillgängligt för dem 24. Såsom
anges i revisionsrättens särskilda rapport nr 28/2018 25 varierar den nivå av stöd som
de nationella kontaktpunkterna erbjuder mellan medlemsstaterna. I vissa länder
arbetar de heltid som nationella kontaktpunkter, medan de i andra måste kombinera
sina uppgifter med andra ansvarsområden.
Evaluation of the SME instrument and the activities under Horizon 2020 Work Programme
Innovation in SMEs, februari 2017.
http://ec.europa.eu/research/participants/data/support/ncp/h2020-standardsprinciples_en.pdf
Särskild rapport nr 28/2018. De flesta förenklingsåtgärder som införts i Horisont 2020 har
gjort livet lättare för stödmottagarna, men det finns fortfarande möjligheter till
förbättringar.
Den nivå av stöd som de nationella kontaktpunkterna erbjuder varierar mellan
medlemsstaterna, vilket påverkar deltagandet och framgångsgraden. I bara två av de
sex medlemsstater som besöktes var de nationella kontaktpunkterna helt fokuserade
på sin roll. De nationella kontaktpunkterna i två medlemsstater anordnade
workshoppar om hur man skriver förslag och förhandsgranskade ansökningar. En
kontaktpunkt lät sökande presentera sina förslag inför en låtsasjury. Andra gjorde inte
mycket förutom att anordna informationsdagar om Horisont 2020.
De nationella kontaktpunkterna och EEN rapporterade att SMF-I i huvudsak hade
marknadsförts på nationell nivå, med begränsat stöd från Europeiska kommissionen,
eftersom programmet inte ger de nationella kontaktpunkterna någon specifik budget
för spridningsinsatser.
Access4SMEs är en åtgärd för samordning och stöd inom Horisont 2020 som ska
underlätta gränsöverskridande samarbete mellan nationella kontaktpunkter för små
och medelstora företag, främja tillgången till riskfinansiering samt uppgradera
kontaktpunkternas kompetens och verktyg så att de kan ge bättre stöd 26.
Intervjuobjekten uppgav att Access4SMEs har varit den främsta källan till information
om SMF-I för de nationella kontaktpunkterna, EEN och stödmottagarna. Nätverket
inrättades dock först i september 2016 – nästan tre år efter det att instrumentet
lanserades – och det existerade alltså inte när dess tjänster hade varit som mest
användbara.
Urval av projekt
Ett ändamålsenligt urvalsförfarande är avgörande för att se till att de bästa
ansökningarna väljs ut för finansiering. Mot denna bakgrund bör urvalsförfarandet ha
tillräckligt med resurser och lämpliga experter utsedda för varje utvärderingssteg.
SMF-instrumentet är baserat på en kontinuerligt öppen förslagsinfordran, med
fyra inlämningsdatum per fas och år. Utvärderingsprocessen utförs på distans av fyra
oberoende utvärderare per förslag. Sedan 2018 har urvalsförfarandet för fas 2-bidrag
inkluderat presentation av projekten för en jury, som ett andra utvärderingssteg som
utförs av en panel bestående av sex experter (investerare för det mesta).
http://www.access4smes.eu/project/#_goal
Begränsade utvärderingsresurser och ett distansutvärderingsförfarande
som är överbelastat på grund av ett stort antal ansökningar
Easme tar emot och handlägger en mängd förslag vid samtliga fyra
inlämningsdatum per år för var och en av de två faserna. Vid det sista
inlämningsdatumet för 2018 tog Easme emot mer än 1 800 ansökningar för fas 2 och
för fas 1.
Utvärderingsprocessen försvåras av en kombination av begränsade resurser och
ett stort antal inlämnade förslag. Utvärderarna har bara 1,6 timmar i fas 1 och
2,4 timmar i fas 2 på sig att slutföra utvärderingen och fylla i tillhörande
dokumentation, trots att ansökningarna är långa (tio sidor exklusive bilagor för fas 1
och 30 sidor exklusive bilagor för fas 2).
I vår enkät svarade bara 34 % av utvärderarna i fas 2 att de 2,4 timmar som
tilldelades av kommissionen för att utvärdera förslagen var tillräckliga. Den
genomsnittliga tid som behövdes var 5,1 timmar. För fas 1 var 56 % av de tillfrågade
nöjda, och det krävdes 3 timmar i stället för de 1,6 timmar som kommissionen
tilldelade (se figur 7).
Figur 7 – Utvärderarnas nöjdhet med antalet timmar som tilldelats för
utvärderingen av förslag
0%
Fas 1
Fas 2
%
%
%
7%
%
%
%
%
%
%
%
%
%
Mycket nöjd
%
%
Nöjd
Inte nöjd
%
9%
%
Inte alls nöjd
Källa: Revisionsrättens enkät till utvärderare.
De utvärderare som svarade på vår enkät var oftast nöjda med den vägledning
och utbildning som erbjöds, men de skulle vilja få återkoppling på sina utvärderingar
och utfallsstatistik, för att lättare kunna riktmärka och förbättra prestationen. De
uttryckte oro kring utbildningen av nya utvärderare och de därav följande
variationerna i poängsättningen. Statistik från Easme bekräftar dessa variationer, och
Horisont 2020-reglerna kräver att 25 % av utvärderarna är nya.
Presentation inför en jury förbättrar i hög grad urvalsförfarandet
samtidigt som tiden för bidragsbeviljande hålls
Införandet av presentationen av projekt för en jury under 2018 var en positiv
förändring. Detta kompenserar för distansutvärderingens inneboende svagheter och
gör det möjligt att verifiera huruvida projektet är praktiskt möjligt och om
arbetsgruppen har potential att genomföra det. Vissa delar är dock fortfarande inte
optimala.
Jurymedlemmarna bedömer 20 projektpresentationer under en
utvärderingsvecka och förväntas läsa de dokument som sökandena lämnar in i förväg.
De jurymedlemmar som intervjuades upplevde dock att de inte fick dokumenten i
tillräckligt god tid för att kunna granska så mycket som 1 600 sidor
ansökningsinformation.
De föreslog också att de skulle få tillgång till kommentarerna i
distansutvärderarnas rapporter. På så sätt skulle användbar kunskap tas tillvara och
effektiviteten förbättras, med tanke på den begränsade tiden för att förbereda och
diskutera projektens jurypresentationer. På liknande sätt ansåg utvärderarna att
kvaliteten på deras utvärderingar skulle förbättras om de fick tillgång till
jurymedlemmarnas kommentarer om de förslag som de hade utvärderat.
Ingen systematisk due diligence-granskning utförs i nuläget av ansökningar som
når presentationsstadiet. Jurymedlemmarna uppgav behovet av en ”lätt” due
diligence-process för att kontrollera om den information som sökandena lämnar om
patent, företagsprofil och arbetsgruppens sammansättning stämmer.
Kommissionen har fastställt målet för tiden för bidragsbeviljande (tiden mellan
inlämningsdatumet och undertecknandet av bidragsavtalet) till högst tre månader för
fas 1 och sex månader för fas 2. Den faktiska tiden för bidragsbeviljandet har minskat
sedan programmet startade, trots införandet av jurypresentationen, och under 2018
undertecknade Easme 90 % av bidragen inom den fastställda tidsperioden.
Vissa it-verktyg utgör en risk för utvärderingsprocessen
De sökande lämnar in förslag online via det elektroniska systemet för inlämning
av förslag på Horisont 2020:s deltagarportal.
För att arrangera projektpresentationer och sätta ihop juryer med lämpliga
färdigheter använder Easme en arbetsbok i ett kalkylprogram, vilken skulle kunna
krascha och därmed orsaka förseningar och äventyra utvärderingsförfarandet.
Eftersom det inte finns något särskilt it-verktyg för att ersätta de sökande för
deras deltagande i presentationen, registreras de som utvärderare i det interna
experthanteringssystemet. Det finns därmed en risk för att de av en händelse
kontaktas för att utvärdera förslag.
Dessutom kräver de ändringar av urvalsprocessen som infördes i september 2019
enligt Europeiska innovationsrådets utökade pilotprojekt (begäran om finansiella
uppgifter från deltagarna och information om teknisk mognadsgrad)
påbyggnadslösningar som fortfarande inte har utvecklats.
Förslag som lämnas in på nytt är betungande för utvärderingsresurserna
Det finns ingen gräns för hur många gånger en icke-utvald ansökan får lämnas in
på nytt till SMF-I. Vid utvärderingen behandlas ett förslag som lämnats in på nytt på
samma sätt som alla andra ursprungliga ansökningar, utan att någon information från
tidigare utvärderingar vidarebefordras.
Den ytterligare kostnad som det innebär för sökanden att lämna in ett oförändrat
förslag är försumbar. Antalet ansökningar som lämnats in på nytt har ökat stadigt och
utgör nu en stor andel av de totala ansökningarna. För de senaste inlämningsdatumen
för fas 2 under 2018 (se figur 8) var 66 % av ansökningarna förslag som lämnades in på
nytt, och hälften av dessa lämnades in för åtminstone tredje gången.
Figur 8 – Antal förslag som lämnas in på nytt i fas 2
%
%
%
%
%
0%
% förslag som skickats in på nytt
% förslag som skickats in minst 3 ggr
Källa: Revisionsrätten, på grundval av uppgifter från kommissionen (fram till slutet av 2018).
Att ansökningarna har ökat med tiden beror bara på att samma förslag lämnas in
igen. Antalet nya projekt som ansöker till fas 2 har legat kvar på 500 ansökningar per
inlämningsdatum (se figur 9).
Figur 9 – Fas 2-projekt: nya jämfört med totalsumman
2 250
2 000
1 750
1 500
1 250
1 000
Totalt antal inlämnade projekt
Nya projekt
Linjär (totalt antal inlämnade projekt)
Linjär (nya projekt)
Källa: Revisionsrätten, på grundval av uppgifter från kommissionen.
Förslag som lämnas in på nytt utgör en betydande och allt större belastning för
utvärderingsresurserna. Mellan 2015 och 2018 var utvärderingskostnaden för förslag
som lämnades in för tredje gången (eller fler) – bara med hänsyn tagen till arvodena
för de expertutvärderare som utför sitt arbete på distans – mer än 4,3 miljoner euro
(inklusive mer än 1,8 miljoner euro under 2018).
Halvtidsutvärderingen av Horisont 2020 tydde på att den överdrivet stora
mängden registrerade ansökningar avskräckte från deltagande, försämrade
utvärderingarnas kvalitet, dränerade resurserna och lämnade ett stort antal
högkvalitativa förslag utan finansiering.
Den genomsnittliga framgångsgraden för inlämnade ansökningar till SMF-I är
4,7 % i fas 2 och 8,6 % i fas 1. Om vi beräknar framgångsgraden per projektförslag
snarare än per inlämning är det dock omkring 11,5 % av fas 2-förslagen och 16,6 % av
fas 1-förslagen som i slutändan väljs ut.
Stödets ändamålsenlighet i SMF-instrumentets faser
Det stöd som beviljas genom SMF-I bör ges i rätt tid, vara relevant och uppfylla
behoven hos innovativa små och medelstora företag.
Fas 1 ger användbart stöd till små och medelstora företag men det finns
redan liknande system i vissa medlemsstater
Enligt olika intressenter som intervjuades har fas 1 och fas 2 i praktiken blivit som
två olika program. Fas 1 hjälper företag som saknar erfarenhet av offentlig finansiering,
till exempel små it-företag eller uppstartsföretag. Fas 2 är mer komplex, vilket innebär
att de företagstyper som ansöker till fas 1 tycker att det är en större utmaning att söka
till fas 2.
Skillnaderna i framgångsgrad mellan företag som går igenom fas 1 innan de
ansöker till fas 2 och företag som ansöker direkt till fas 2 har jämnats ut under
genomförandet av SMF-I. Men framgångsgraden för fas 2 är fortfarande 50 % högre
för företag som går igenom fas 1 än för företag som ansöker direkt till fas 2 (se
figur 10).
Figur 10 – Jämförelse av framgångsgraden för små och medelstora
företag som ansöker direkt till fas 2 och små och medelstora företag som
redan har ansökt till fas 1 innan fas 2
9%
8,41 %
7,68 %
8%
7%
5,97 %
6%
5%
4%
3%
2%
5,32 %
5,04 %
4,05 %
3,94 %
3,93 %
3,13 %
5,12 %
4,28 %
3,68 %
3,74 %
2,88 %
2,87 %
1%
0%
Framgångsgrad direkt inlämning
Framgångsgrad efter fas 1
Framgångsgrad sammantaget
Källa: Revisionsrätten på grundval av uppgifter från Easme.
Fas 2-mottagare som hade gått igenom genom fas 1 uppgav att den första fasen
var en bra förberedelse, som hjälpte dem att förbättra projektet.
I vissa medlemsstater ansåg intressenter som intervjuades att fas 1-projekt ofta
hade kunnat utföras lika väl på nationell nivå, även om detta skulle vara en utmaning i
vissa medlemsstater.
I vår enkät till de nationella innovationsmyndigheterna uppgav 48 % av de som
svarade att deras medlemsstat hade nationella program som liknade fas 1. När vi
frågade dem om de främsta styrkorna hos den första fasen av SMF-I jämfört med de
nationella programmen uppgav myndigheterna snabba och öppna urvalsförfaranden,
den trovärdighet som EU:s varumärke medför och tillgången till coachning och
företagsacceleration. Dessutom lovordade de den kritiska massa av innovativa företag
som hade skapats tack vare den första fasen av SMF-I, som hade lyckats locka till sig
många innovativa företag till EU-programmet.
När vi bad om deras synpunkter på huruvida fas 1 borde fortsätta under det nya
ramprogrammet svarade 86 % av de nationella innovationsmyndigheterna att fas 1
borde behållas under det nya ramprogrammet (se ruta 1 för exempel på nationella
innovationsmyndigheters åsikter om huruvida man borde fortsätta att finansiera
fas 1). De som ställde sig positiva till att fas 1 skulle fortsätta uppgav att
företagsaccelerations- och coachningstjänsterna hade förbättrat dessa företags
kapacitet att hantera innovationsverksamhet på ett professionellt sätt och gjort det
möjligt för dem att skala upp och växa. De menade att förslagsinfordrans europeiska
karaktär sporrade små och medelstora företag att höja sin ambitionsnivå från de
inledande utvecklingsstadierna, och att den enkla och snabba utvärderingsprocessen
saknade motsvarigheter på nationell nivå. De som var emot att fas 1 skulle fortsätta
(14 %) noterade att den inte hade något mervärde jämfört med nationella/regionala
instrument och att det inte fanns någon påtaglig koppling mellan fas 1 och fas 2.
Ruta 1
De nationella innovationsmyndigheternas åsikter om fas 1
—
Fas 1 har varit en utmärkt inkörsport till Horisont 2020 för små och
medelstora företag som saknat erfarenhet från europeiska eller
internationella forsknings- och innovationsprogram. De
företagsaccelerations- och coachningstjänster som EEN tillhandahållit små
och medelstora företag har förbättrat företagens kapacitet att hantera
innovationsverksamhet på ett professionellt sätt och gjort det möjligt för
dem att skala upp och växa.”
—
Fas 1 har gjort det möjligt för små och medelstora företag att utvecklas.
Sådana företag saknar ofta kunskap och resurser att göra omfattande
undersökningar av immaterialrättigheter, marknader och konkurrens och så
vidare. När de har slutfört fas 1-projektet är de också väl förberedda att inte
bara ansöka om fas 2-finansiering, utan även skaffa andra
finansieringsresurser/annat kapital. Det bidrag som erhålls från
kommissionen är också en slags pålitlighets- och kvalitetsstämpel.”
—
Fas 1 är värdefull men gör inte mest nytta. Det är snarare viktigt att
medlemsstaterna/de associerade länderna också investerar själva, så att
småskaliga insatser som denna kan lämnas till de nationella/regionala
myndigheterna. Alla medlemsstater har dock inte möjlighet att ge sådant
stöd.”
—
Fas 1 ger ingen additionalitet – alla medlemsstater kan inrätta ett liknande
program.”
Fas 1 är alltför betungande för förvaltningen av SMF-instrumentet
Sedan SMF-I inleddes har 3 978 fas 1-bidragsavtal undertecknats. Arbetet från
start till slut kräver avsevärda administrativa insatser i form av utvärdering,
bidragsförberedelser, undertecknande av bidrag och coachningstjänster. Fyra
projekthandläggare har hand om omkring 1 000 projekt om året. Projektövervakningen
är därför begränsad till administrativa kontroller och man bedömer alltså inte
genomförbarhetsstudiens kvalitet.
Tabell 1 jämför vad distansutvärderingen kostar per fas med de sammanlagda
belopp som beviljats. Där framgår att det är stor skillnad mellan kostnaderna för de
olika faserna, då de relativa utvärderingskostnaderna är tio gånger högre (per beviljad
euro) i fas 1 än i fas 2. Riktmärket för utvärderingskostnaden inom sektorn för privat
riskkapital är 3 %.
Tabell 1 – Kostnad för distansutvärderingar
FAS 1
FAS 2
EUR
EUR
Total kostnad
840 EUR
200 EUR
Beviljat belopp
000 EUR
609 479 EUR
8,3 %
0,7 %
Antal utvärderade förslag
Antal utvärderade förslag per dag och utvärderare
Kostnad för distansutvärdering per förslag
Utvärderingskostnad/beviljat belopp
Källa: Revisionsrätten.
Trots de större administrativa omkostnaderna i fas 1 jämfört med fas 2
tillhandahåller fas 1 ändamålsenligt stöd tack vare den snabba urvalsprocessen på EUnivå, EU-varumärket för stödmottagarna och tillgången till
företagsaccelerationstjänsterna. Dessutom har den lockat till sig många innovativa
företag till EU-programmet. I länder där det redan finns program som liknar fas 1
minskar instrumentets relevans.
Kommissionen har lagt ner fas 1 från och med september 2019.
Fas 2 ger ändamålsenligt stöd till små och medelstora företag
De intressenter som intervjuades (representanter från nationella
innovationsmyndigheter och nationella kontaktpunkter, innovationsexperter,
utvärderare, jurymedlemmar, EEN, paraplyorganisationer för små och medelstora
företag och stödmottagare) var eniga i sitt gillande av fas 2 på grund av de många
positiva inslagen, till exempel följande:
—
Stora ekonomiska stöd vid en hög teknisk mognadsgrad som medlemsstaterna
inte kan ge 27.
—
Konkurrensen bland små och medelstora företag på EU-nivå.
—
Möjligheten att locka till sig ytterligare investeringar med hjälp av EU-varumärket
(se punkterna 119 och 121).
—
Tillgången till coachning och tjänster för företagsacceleration.
—
Enkla och snabba urvals- och tilldelningsprocesser jämfört med de nationella
systemen.
—
Fokus på projektens marknadslanseringsstrategi, där man tar fram en
handlingsplan som specificerar hur företaget ska nå kunderna och uppnå en
konkurrensmässig fördel.
I vår enkät till de nationella innovationsmyndigheterna frågade vi dem huruvida
de tyckte att den andra fasen av SMF-I borde fortsätta inom ramen för
Horisont Europa och varför (se ruta 2 för exempel på dessa myndigheters synpunkter
på huruvida man borde fortsätta att finansiera fas 2). Alla svarande sa att den borde
fortsätta.
Kommissionens förordning (EU) nr 651/2014 genom vilken vissa kategorier av stöd förklaras
förenliga med den inre marknaden.
Ruta 2
De nationella innovationsmyndigheternas åsikter om fas 2
—
Fas 2 erbjuder något som skiljer sig från vad som finns tillgängligt på nationell
nivå. Den underlättar också skapandet av internationella nätverk. Det är
också viktigt med coachning.
—
Fas 2 är ett mycket bra instrument som är lätt för sökandena att förstå.
—
Fas 2 är ett viktigt och unikt program när det gäller att stödja växande små
och medelstora företag under pilotfasen.
—
Systemets framgång och popularitet bland små och medelstora företag har
bevisat att det har en mycket lämplig struktur för dessa företag. De
förändringar som gjordes under genomförandeperioden (i synnerhet
intervjuer) har höjt systemets värde.
När myndigheterna rådfrågades om huruvida man borde förändra utformningen
av SMF-I avsevärt svarade 75 % ”nej”, 16 % tyckte att det räckte med begränsade
förändringar och bara 11 % menade att mer djupgående förändringar krävdes. Detta
tyder på att den nuvarande form som fas 2 har i allmänhet är väl uppskattad.
Fas 2 av SMF-I ger ändamålsenligt stöd till stödmottagarna. Den ger projekten
EU:s varumärke, vilket innebär synlighet för företagen och projekten, hjälper dem att
anskaffa ytterligare investeringar och ger tillgång till EU-nätverket för coachning och
företagsaccelerationstjänster. Fas 2 uppskattas stort i sin nuvarande form bland de
nationella innovationsmyndigheter som deltog i enkäten. Denna åsikt delades av alla
intressenter som intervjuades.
Företagsaccelerationstjänsterna i fas 3 har potential, men de lanserades
sent
Coachningen och företagsaccelerationstjänsterna (fas 3) spelar en viktig roll i
SMF-instrumentets övergripande struktur eftersom de syftar till att uppfylla de små
och medelstora företagens innovationsbehov genom skräddarsytt stöd,
kompetensutveckling och arbete i nätverk. Enligt en studie som offentliggjorts av
University of Manchester lyckas företag (särskilt små företag) mycket bättre via
åtgärder som kombinerar direkt och indirekt stöd 28.
Coachningen omfattar en rad olika ämnen, framför allt affärsutveckling,
organisationsutveckling, samarbete och finansiering. Stödmottagarna i fas 1 fick tre
dagars coachning och stödmottagarna i fas 2 fick tolv. SMF-I har lett till att man
inrättat det första europeiska nätverket av coacher för att stödja stödmottagarna.
Företagsaccelerationstjänsterna är öppna för både fas 1- och fas 2-stödmottagare
och inbegriper deltagande i följande tjänster:
—
Mässor och konferenser.
—
Företagsdagar.
—
Evenemang för investerare.
—
Toppmötet EIC Innovators.
—
Mentorskap.
—
Samverkansplattformen för EIC.
—
Ett verktyg för matchning med investerare.
—
EIC Academy.
The Impact of Direct Support to R&D and Innovation in Firms”, Compendium of Evidence
on the Effectiveness of Innovation Policy Intervention, augusti 2012.
Evenemang och andra företagsaccelerationstjänster i fas 3 har främst fokuserat
på att skapa förbindelser mellan små och medelstora företag och potentiella
investerare eller affärspartner. Easme har inte gjort särskilt mycket för att hjälpa
stödmottagarna att nå ut till potentiella kunder (såsom stora privata företag eller
offentliga organ genom innovativ offentlig upphandling).
De stödmottagare (små och medelstora företag) som svarade på vår enkät
uppskattade i hög grad både coachningssystemet och alla
företagsaccelerationstjänster som de hade använt (se figur 11). Denna positiva åsikt
bekräftades av våra besök hos stödmottagare och av de nationella
innovationsmyndigheter som deltog i enkäten. De nationella
innovationsmyndigheterna och EEN-knutpunkterna föreslog ändå att Easme skulle
kunna
—
samordna anordnandet av evenemang med lokala aktörer (nationella
innovationsmyndigheter och EEN-knutpunkter) på ett bättre sätt,
—
rikta marknadsföringen av företagsaccelerationstjänsterna bättre för att undvika
att mejla små och medelstora företag om evenemang som inte är relevanta för
dem,
—
utforska möjligheterna att samarbeta med nationella investeringsbanker som
skulle kunna erbjuda SMF-I-stödmottagarna investeringsmöjligheter.
Figur 11 – Stödmottagarnas nöjdhet med coachningen och
företagsaccelerationstjänsterna
0%
%
%
%
%
%
Företagscoachning
Evenemang för investerare
Företagsdagar
Mässor
och konferenser
Toppmötet
EIC Innovators
Verktyg
för matchning med investerare
Samverkansplattformen
för EIC
EIC Academy
Mycket användbar
Användbar
Lite användbar
Inte användbar
Källa: Revisionsrättens enkät till stödmottagare.
De innovationsexperter som intervjuades anser att
företagsaccelerationstjänsterna borde stimulera efterfrågesidan genom att matcha
små och medelstora företag med potentiella stora företagskunder och stödja deras
deltagande i innovativa offentliga upphandlingssystem.
Som en jämförelse är fas 3 av SBIR-programmet inriktat på offentlig
upphandling. I USA måste federala myndigheter med årliga FoU-budgetar som
överskrider 100 miljoner US-dollar anslå 3,2 % till stödmottagarna inom ramen för
SBIR-programmet genom offentlig upphandling. Under 2015 uppgick de kontrakt som
undertecknades mellan federala myndigheter i USA och SBIR-stödmottagarna till
1,3 miljarder US-dollar, medan bidragen sammantaget var värda 1,2 miljarder USdollar 29.
SBA Office of Investment & Innovation om SBIR, december 2016.
Den betydelse som offentlig upphandling har för små och medelstora företag
och uppstartsföretag erkänns av kommissionen i dess vägledning om
innovationsupphandling 30. I detta dokument anges det att ”[g]enom att agera som
banbrytande konsumenter kan offentliga upphandlare ge innovativa företag möjlighet
att testa sina nya lösningar under verkliga förhållanden. Genom att bli deras kunder
och därmed öka deras omsättning kan upphandlande myndigheter dessutom
uppmuntra andra investerare – såväl offentliga som privata – att investera i deras
verksamhet”. I nuläget har dock kommissionen inte inkluderat några system för
innovativ offentlig upphandling bland företagsaccelerationstjänsterna för att skapa
kopplingar mellan SMF-I:s stödmottagare och EU-byråer eller nationella institutioner.
Utnyttjandet av de olika företagsaccelerationstjänsterna har varit lågt. Av de
stödmottagare som ingick i undersökningen deltog 12 % i EIC Academy och 40 % vid
mässor och konferenser (se figur 12). Detta förklaras delvis med att vissa tjänster
startades först i slutet av 2017, nästan fyra år efter det att instrumentet lanserades.
Kommissionens tillkännagivande C(2018) 3051, 15.5.2018.
Figur 12 – Procentandel svarande som inte utnyttjade
företagsaccelerationstjänsterna
EIC Academy
Verktyg för matchning med investerare
Samverkansplattformen för EIC
Evenemang för investerare
Toppmötet EIC Innovators
Företagsdagar
Mentorskap
Mässor & konferenser
% 10 % 20 % 30 % 40 % 50 % 60 % 70 % 80 % 90 % 100 %
Källa: Revisionsrättens enkät till stödmottagare.
SMF-instrumentets ändamålsenlighet har inte bedömts, och dess
framtida roll i Horisont Europa har ännu inte fastställts
För att kunna lämna bidrag i rätt tid till utarbetandet av den nya förordningen
utförde kommissionen flera utvärderingar under SMF-I:s första år – trots att det
saknades mogna uppgifter (se figur 13) – såsom följande:
—
Den halvtidsutvärdering av SMF-I som offentliggjordes i februari 2017, då ännu
inga innovationsprojekt i fas 2 hade slutförts.
—
Den halvtidsutvärdering av Horisont 2020 som offentliggjordes i maj 2017, som
påverkades av samma tidsmässiga begränsningar som i punkten ovan.
—
Den konsekvensbedömning av Horisont Europa som offentliggjordes i juni 2018.
Bara omkring 200 företag hade vid denna tidpunkt slutfört sina
innovationsprojekt i fas 2. Dessutom tar det normalt sett några år att se ett
innovationsprojekts verkliga effekter.
Figur 13 – Samlat antal projekt i SMF-I fas 2 som slutförts och den period
som omfattas av utvärderingen
Uppskattade siffror
1 400
1 200
1 000
Konsekvensbedömning av Horisont Europa
Halvtidsutvärdering av Horisont 2020
Utvärdering av SMF-I
Källa: Revisionsrätten, på grundval av uppgifter från kommissionen.
Eftersom programmet är nytt och det saknas tidigare resultatuppgifter
utvärderades SMF-I endast på grundval av indata och slutförda fas 1-projekt, och inte
på grundval av resultat från fas 2-projekt. De samråd som hölls och de oberoende
rapporter som togs fram för utformningen av Europeiska innovationsrådet inom ramen
för Horisont Europa (se bilaga II) omfattades av samma begränsningar. Därför kunde
kommissionen inte basera utformningen av Europeiska innovationsrådet inom
Horisont Europa på en övergripande analys av SMF-I:s genomförande, uppnådda
resultat och effekter.
Locka till sig investeringar efter finansieringen genom SMFinstrumentet
Ett av syftena med SMF-I är att underlätta tillgången till privat kapital och att
skapa länkar till EU-stödda finansieringsinstrument 31. Enligt rådets beslut 2013/743/EU
planeras ”[l]änkar till finansiella instrument  till exempel genom att prioritera små
och medelstora företag som framgångsrikt har slutfört fas 1 och/eller 2 inom en
öronmärkt volym av finansieringsresurserna”.
Förordning (EU) nr 1291/2013 om inrättande av Horisont 2020.
Kommissionen har bara begränsad kunskap om stödmottagarnas
övergripande finansieringsbehov och har inte skapat länkar till EU:s
finansieringsinstrument
Easme samlar inte systematiskt in information om fas 2-stödmottagarnas
ytterligare finansiella behov för att de ska kunna utveckla sina projekt fullt ut. Easme
utförde under 2016 en enkätundersökning för att bedöma behoven, men ställde inga
frågor om vilken källa som föredrogs eller om hur finansieringen skulle användas.
År 2018 bad GD Forskning och innovation EIB att ta fram en studie om
tillgången till finanser för SMF-I-stödmottagare, som sedan användes för
konsekvensbedömningen av Horisont Europa 32. EIB baserade rapporten på
förhandsbedömningar och på en enkätundersökning bland ett urval av stödmottagare.
Urvalet var dock inte representativt och det vara bara 24 stödmottagare som svarade
på enkäten. Därmed ger rapporten bara begränsad insyn i de faktiska finansiella
behoven hos SMF-I:s stödmottagare.
Vår representativa enkät (se bilaga I) gav en fingervisning om vad fas 2stödmottagarna har för finansiella behov. Framför allt konstaterades följande:
—
Tre fjärdedelar av de som svarade sa att de behövde ytterligare finansiering på i
genomsnitt 7,1 miljoner euro.
—
% av de som svarade som sökte ytterligare finansiering uttryckte intresse för
privata riskkapitalinvesteringar, medan 48 % var öppna för skuldinstrument som
lån eller kreditlinor.
De finansieringsslag som söktes varierar enligt företagsmognad, där unga små
och medelstora företag är mer intresserade av kapitaltillskott än äldre (se figur 14).
Den rådgivande gruppen för EIB-Innovfin: Improving Access to Finance for Beneficiaries of
the SME Instrument, mars 2018.
Figur 14 – Andel svarande som söker stöd i form av riskkapital efter
företagets ålder
0%
< 5 år
5–9 år
10–19 år
≥ 20 år
%
%
%
%
%
Nej
Ja
Källa: Revisionsrättens enkät till stödmottagare.
Majoriteten av SMF-I:s stödmottagare skulle behöva ytterligare finansiering för
att stödja sitt innovationsarbete och lansera sina innovationsprojekt på marknaden.
Kommissionen har dock begränsad kunskap om stödmottagarnas finansiella behov.
Under den fleråriga budgetramen för 2014–2020 lanserade EU ett stort antal
finansieringsinstrument för att stödja innovation i små och medelstora företag33. 64 %
av de stödmottagare som svarade på enkäten kände dock inte till dessa instrument.
Bland annat initiativet för tillgång till riskfinansiering (InnovFin) inom ramen för
Horisont 2020, tillgång till finansiering för små och medelstora företag (Cosme) och
Europeiska fonden för strategiska investeringar (Efsi).
I EIB:s rapport om tillgång till finansiering för SMF-I:s stödmottagare34 drogs
följande slutsatser, som bekräftades genom vår enkät till och intervjuer med
stödmottagare:
—
Det finns ett likviditetsgap för SMF-I-stödmottagarna när projekten lämnar fas 2.
—
Bidragen ger en positiv marknadssignal till privata kapitalgivare.
—
Den tillgängliga informationen om finansieringsinstrument är splittrad och
kommunikationen mellan privata och offentliga kapitalgivare är begränsad.
En EAG-rapport35 från 2016 framhöll bristen på synergier mellan EU:s olika
finansiella insatser och behovet av att samordna SMF-I med andra offentliga
investerare för att bättre kunna bemöta projektens förfrågningar om medel när fas 2
hade slutförts.
Vi analyserade den förteckning över mottagare av riskkapital med EU-stöd som
sammanställs av EIB och EIF och konstaterade att i slutet av 2018 hade bara 16 SMF-Istödmottagare (varav åtta befann sig i fas 2) fått sådant ekonomiskt stöd. I fem fall
gjordes finansieringsinstrumentets investering innan bidraget från SMF-I hade
beviljats.
Ett av målen med SMF-I har sedan start varit att skapa länkar till EU-stödda
finansieringsinstrument. Kommissionen har dock gjort mycket lite för att uppnå detta:
den öronmärkte inte några medel för SMF-I-stödmottagarna, och stödmottagarna har
begränsad kännedom om EU-stödda finansieringsinstrument.
Den rådgivande gruppen för EIB-Innovfin: Improving Access to Finance for Beneficiaries of
the SME Instrument, mars 2018.
H2020 EAG, Innovation in SMEs, Annual Report 2016.
Stödmottagarna lockar till sig ytterligare investeringar, men nivåerna
varierar i EU
De bidragsavtal som tecknas via SMF-I kräver inte att stödmottagarna
rapporterar när väl projektet har slutförts. Easme övervakar i stället hur
stödmottagarna utvecklas efter det att SMF-I-bidraget tilldelades genom två
databaskällor, som sköts av externa uppdragstagare:
—
Källa 1 används för att bedöma de investeringar som SMF-I-stödmottagarna har
anskaffat. Databasen sammanställs genom insamling av information om
investeringsrundor som finns offentligt tillgänglig online. För att bedöma hur pass
tillförlitlig denna källa är kontrollerade vi ett slumpmässigt urval på 30 fas 2stödmottagare, vilket bekräftade siffrorna från den tillgängliga informationen
online.
—
Källa 2 används för att bedöma utvecklingen över tid av SMF-I-stödmottagarnas
prestation i fråga om omsättning, nettointäkter, kassaflöde och
sysselsättningsnivåer.
Information som samlas in direkt från stödmottagarna kan vara mindre
tillförlitlig då självrapporteringen kan vara vinklad. Dessutom är användningen av
tredjepartsinformation mer kostnadseffektiv. Samtidigt är dock båda dessa
informationskällor ofullständiga eftersom
—
källa 1 underskattar de faktiska investeringar som SMF-I-stödmottagarna har
anskaffat, eftersom man inte vet hur mycket investeringar i form av skulder och
kapitaltillskott (som inte offentliggörs online) som har anskaffats,
—
källa 2 tillhandahåller fullständiga uppgifter för bara omkring 60 % av alla SMF-Istödmottagare 36.
Enligt den information som finns tillgänglig online är förhållandet mellan
investeringar och bidrag 2,9 för fas 2-stödmottagare som fick bidrag från SMF-I under
och 2015 och som slutförde sina innovationsprojekt 2017. Figur 15 visar
utvecklingen i fråga om de ytterligare investeringar som stödmottagarna anskaffat
under åren efter det att SMF-I-stödet beviljades.
Källa: Easme.
Figur 15 – Utveckling i fråga om de ytterligare investeringar som
stödmottagarna anskaffat under åren efter bidraget
1 000
Miljoner euro
1 år
2 år
3 år
4 år
5 år
-
Källa: Revisionsrätten på grundval av uppgifter från Easme.
Dessa siffror inkluderar inte investeringsrundor som inte publiceras online,
såsom majoriteten av alla mindre kapitaltillskott och nästan allt skuldkapital som
tillhandahålls av banker, fonder och andra finansiella aktörer. Uppgifter om anskaffade
investeringar finns offentligt tillgängliga online för bara 11 % av alla fas 2stödmottagare.
Jämförelsevis uppgav majoriteten av alla fas 2-stödmottagare (78 % av de som
svarade på vår enkät) att fas 2-finansieringen hade hjälp dem att mobilisera ytterligare
finansiering för att stödja deras innovationsbehov. Stödmottagarnas faktiska förmåga
att locka till sig investeringar är därför antagligen större än vad som framgår av den
information som finns tillgänglig online.
Enligt information från en tredje part (källa 1, se punkt 117) som bekräftades
genom uppgifter som samlades in i samband med projektrapporteringen uppvisar
SMF-I-stödmottagarna positiva tendenser i fråga om strukturell tillväxt. Omkring 75 %
av företagen hade upplevt en ökning av sina rörelseintäkter sedan de ansökte om
bidraget, och 67 % hade ökat sin personalstyrka.
En gedigen uppsättning effektmått som baseras på tillförlitliga uppgifter,
kombinerat med helt automatisk profilering av de företag som lämnar in projektförslag
och väljs ut för bidrag, är nödvändig för att utveckla en ändamålsenlig
affärsunderrättelsestrategi. Detta skulle kunna hjälpa till med följande:
—
Fastställa mönster för deltagande och potentiella obalanser.
—
Koppla effektmått till deltagarkluster genom att tillhandahålla värdefull
information om hur instrumentets övergripande effekter kan maximeras.
SMF-I har under det utökade pilotprojektet för ett europeiskt innovationsråd
förbättrat företagsprofileringen eftersom de nya administrativa formulären samlar in
uppgifter om tidigare investeringsrundor, finansiella uppgifter och ägarstrukturen hos
de som lämnar förslagen. Hittills har man dock inte systematiskt samlat in information
om aktieägarnas kön i det skede då förslagen lämnas in, vilket är ett av de kriterier som
bedöms av jurymedlemmarna.
Det finns betydande skillnader mellan de deltagande länderna, där fas 2-
deltagarna i nordvästra Europa lyckas anskaffa mer privata resurser än små och
medelstora företag i södra och östra Europa (se figur 16)37. Dessa obalanser kan delvis
förklaras med skillnaderna mellan riskkapitalmarknaderna i dessa länder.
Källa: Revisionsrätten baserat på uppgifter från Easme. Länder för vilka inga ytterligare
investeringar har kunnat konstateras genom webbsökningar har inte tagits med i tabellen.
Figur 16 – Genomsnittliga investeringar som anskaffats per fas 2stödmottagare, per mottagarland
(I miljoner euro)
Finland
Nederländerna
Tyskland
Förenade kungariket
Estland
Sverige
Israel
Irland
Frankrike
Island
Spanien
Portugal
Norge
Danmark
Italien
Belgien
Polen
Källa: Revisionsrätten på grundval av uppgifter från Easme.
Resultatet av vår enkät till stödmottagarna tyder på att den geografiska platsen
är en avgörande faktor som påverkar hur pass benäget ett företag är att söka efter
kapital- och/eller skuldinvesteringar. I de nordiska länderna och i Förenade kungariket
planerade 84 % av alla tillfrågade att söka efter kapitaltillskott, jämfört med 54 % i
Spanien och 42 % i Italien.
EAG:s rapport om SMF-I tog upp frågan om variationer mellan länder och olika
kulturer vad gäller användningen av marknadsbaserade instrument, och
rekommenderade en kartläggning av det europeiska landskapet för att få mer kunskap
om potentiella medinvesterare och för att kontrollera om gränsöverskridande aktörer
kan överbrygga vissa finansieringsunderskott när de nationella systemen inte fungerar.
Plattformar och särskilda evenemang skulle kunna hjälpa till med denna process 38.
Bild 3 visar flödet av ytterligare investeringar över 10 miljoner euro till
stödmottagande länder, uppdelat efter ursprungsland. Av de 1,8 miljarder euro i
ytterligare investeringar som fas 2-stödmottagarna har anskaffat (se punkt 119)
kommer cirka 400 miljoner euro från investerare med säte i USA och 181 miljoner euro
från investerare i Kina. Den största enskilda investeraren i fas 2-stödmottagare har sitt
säte i USA, och tre av de fem största investeringarna (över 50 miljoner euro) kommer
från investerare utanför EU.
H2020 EAG, Innovation in SMEs, Consultation on the EU Strategic WP 2018–2020, juni 2016.
Bild 3 – Investeringar som anskaffats per investerarland och
stödmottagarland i miljoner euro
INVESTERARE
STÖDMOTTAGARE
Finland
USA
403,0
391,0
Förenade kungariket
206,1
Tyskland
330,6
Nederländerna
198,5
Förenade kungariket
Kina
252,3
180,9
Sverige
104,1
Nederländerna
Frankrike
241,3
87,2
Okänt
75,1
Sverige
116,0
Hongkong
74,4
Israel
81,9
Finland
68,9
Irland
Tyskland
62,0
64,2
Frankrike
Luxemburg
58,0
41,7
Israel
33,4
Spanien
Spanien
25,2
Estland
Andra*
Norge
51,8
15,0
12,5
73,6
*
Norge
Schweiz
Irland
Belgien
Sydafrika
Japan
15,3
14,7
12,0
10,9
10,7
10,0
» Sverige
» Tyskland
» Irland
» Nederländerna
» Förenade kungariket
» Spanien
Källa: Revisionsrätten på grundval av uppgifter från Easme.
EU
Associerade länder till
Horisont 2020
Övriga länder
Slutsatser och rekommendationer
Vi konstaterade att SMF-instrumentet ger ändamålsenligt stöd till små och
medelstora företag när de utvecklar sina innovationsprojekt. EU:s varumärke hjälper
dessutom företagen att locka till sig ytterligare investeringar. Det har dock inte skapats
länkar till EU-stödda finansieringsinstrument som skulle kunna hjälpa stödmottagarna
att skala upp och lansera sina innovationsprojekt på marknaden. Både fas 1 och fas 2
av instrumentet ger små och medelstora företag ändamålsenligt stöd, men fas 1
medför oproportionerligt höga administrativa kostnader. Instrumentet förvaltas av
kommissionen på ett kompetent sätt. Det stora antal ansökningar som lämnas in på
nytt och de begränsade resurserna har hindrat urvalsförfarandet och utvecklingen av
företagsaccelerationstjänsterna.
Alla rekommendationer är tillämpliga på efterträdaren till SMF-instrumentet
inom ramen för Horisont Europa.
Inriktning på rätt stödmottagare
Instrumentets breda syften och mål har, tillsammans med de ändringar som
gjorts under dess genomförande, skapat ovisshet bland berörda parter. Den nuvarande
företagsprofilen passar den akademiska modellen med företag med tillväxtpotential,
men instrumentet finansierar vissa små och medelstora företag som skulle kunna ha
finansierats av marknaden (se punkterna 28–39).
Geografisk täckning
Deltagandet i instrumentet varierar påtagligt mellan länderna, delvis på grund
av faktorer som kommissionen inte kan kontrollera, men också på grund av de
varierande nivåerna av stöd från de nationella kontaktpunkterna och Enterprise
Europe Network (se punkterna 43 och 45 och figur 5). Med en begränsad budget
organiserade kommissionen evenemang och kommunikationsverksamheter, men dess
marknadsföring och kommunikation var varken strukturerad eller tillräckligt välriktad
för att nå rätt företag (se punkterna 40–58).
Rekommendation 1 – Förbättra kommunikationsstrategin och
stödet till de nationella kontaktpunkterna, i synnerhet för de
medlemsstater som har lägst deltagande
Kommissionen bör
fokusera mer på en marknadsförings- och kommunikationsstrategi för att öka
medvetenheten bland de små och medelstora företag som utgör målgruppen om
de finansieringsmöjligheter som erbjuds av instrumentet och dess efterträdare
under Horisont Europa,
förbättra sitt stöd till de små och medelstora företagens nationella
kontaktpunkter och till Enterprise Europe Network genom att främja projekt för
ömsesidigt lärande och utbyten av bästa praxis och säkerställa att stödet till de
nationella kontaktpunkterna för små och medelstora företag är på plats när nästa
ramprogram inleds.
Måldatum för genomförande: 2021
Urval av projekt
Utvärderings- och urvalsförfarandena har förbättrats under instrumentets
livstid. Presentationen inför en jury har varit särskilt nyttig när det gäller att identifiera
de bästa förslagen samtidigt som man håller tidsmålet för beviljande av bidrag (se
punkterna 65–69).
Det förekommer variationer i de poäng som tilldelas i distansutvärderingarna,
vilket delvis kan förklaras med de begränsade resurserna och det stora antalet förslag
som lämnas in. Utbildningen för utvärderarna uppskattas mycket, men ytterligare
återkoppling efterfrågas på olika nivåer. De it-verktyg som används är inte lämpade för
ändamålet och äventyrar utvärderingsprocessen (se punkterna 61–64 och 70–73).
Att förslag som inte blivit godkända lämnas in på nytt utgör en stor och ökande
belastning för förvaltnings- och utvärderingsresurserna och ökar de administrativa
kostnaderna. Dessutom sänker detta framgångsgraden, det vill säga andelen
ansökningar som beviljas stöd, vilket i sin tur avskräcker från deltagande (se
punkterna 74–79).
Rekommendation 2 – Förbättra urvalsförfarandet
För att optimera resursanvändningen och säkerställa ett effektivt urval av de bästa
förslagen bör kommissionen förbättra urvalsförfarandet på följande sätt:
Ge distansutvärderarna mer tid för att utföra sitt arbete.
Inrätta en tvåvägskanal för information mellan distansutvärderarna och
jurymedlemmarna för att låta de sistnämnda få tillgång till distansutvärderingen
och ge de förstnämnda återkoppling om kvaliteten på deras arbete.
Utveckla skräddarsydda it-verktyg för att kunna sköta utvärderingsprocessen på
ett tillförlitligt sätt.
Begränsa antalet gånger ett förslag får lämnas in på nytt, för att på så sätt frigöra
resurser som i nuläget används för att utvärdera samma förslag på nytt vid flera
på varandra följande inlämningsdatum.
För att uppmuntra fler små och medelstora företag med utmärkta
innovationsprojekt att delta borde kommissionen offentliggöra framgångsgraden
per projektförslag.
Måldatum för genomförande: 2021
Stödets ändamålsenlighet i SMF-instrumentets faser
Fas 1 ger ändamålsenligt stöd, tack vare den snabba urvalsprocessen, EU:s
varumärke för stödmottagarna och tillgången till företagsaccelerationstjänster.
Dessutom har den lockat till sig många innovativa företag till EU-programmet. Den
innebär dock en överdriven börda för kommissionens förvaltning av instrumentet och
det finns länder som redan har liknande program (se punkterna 81–89). Fas 1 avbröts
från och med september 2019.
Fas 2 av SMF-I ger ändamålsenligt stöd till stödmottagarna och är mycket
uppskattad bland alla intressenter i sin nuvarande form. Den ger projekten EU:s
varumärke, vilket innebär synlighet för företagen och projekten, hjälper dem att
anskaffa ytterligare investeringar och ger tillgång till EU-nätverket av coachning och
företagsaccelerationstjänster (se punkterna 91–94).
Rekommendation 3 – Ersätt fas 1 och bygg vidare på fas 2stödet till små och medelstora företag
Kommissionen bör
föreslå för medlemsstaterna att kommissionen ska förvalta ett system som liknar
fas 1,
ge stödmottagarna i det systemet tillgång till coachning och
företagsaccelerationstjänster samt EU:s varumärke,
bevara ett system som liknar fas 2 inom Europeiska innovationsrådet inom ramen
för Horisont Europa, och bygga vidare på resultaten från
Europeiska innovationsrådets pilotprojekt.
Måldatum för genomförande: 2021
Tjänsterna för coachning och företagsacceleration kan förstärka instrumentets
effekter men de lanserade sent, är inte tillräckligt synliga och det var bara en liten
andel av de små och medelstora företagen som använde sig av tjänsterna. De tilldelade
resurserna är begränsade och tjänsterna skulle kunna vara mer skräddarsydda och
bättre riktade mot efterfrågesidan (se punkterna 95–103).
Rekommendation 4 – Förbättra företagsaccelerationstjänsterna
Kommissionen bör förbättra företagsaccelerationstjänsterna genom att anslå lämpliga
resurser till detta område, för att
tillhandahålla mer skräddarsydda företagsaccelerationstjänster,
öka medvetenheten bland stödmottagarna med hjälp av en riktad
kommunikationsstrategi,
hantera efterfrågesidan på ett bättre sätt genom att etablera kontakt med stora
privata kunder och genom offentlig upphandling för innovativa projekt.
Måldatum för genomförande: 2022
Locka till sig investeringar efter finansieringen genom SMF-instrumentet
Majoriteten av stödmottagarna behöver fortfarande ytterligare finansiering för
att stödja sitt innovationsarbete och lansera sina innovationsprojekt på marknaden.
Kommissionen har dock inte gjort mycket för att skapa länkar till EU-stödda
finansieringsinstrument och har inte utforskat samarbetsmöjligheter med nationella
investeringsbanker. Dessutom är stödmottagarna ofta omedvetna om de EU-stödda
finansieringsinstrument som finns, och kommissionens kunskap om stödmottagarnas
finansiella behov är begränsad. EIB:s rapport från 2018 om tillgång till finansiering för
stödmottagare bekräftade att den tillgängliga informationen om
finansieringsinstrument är splittrad och att kommunikationen mellan privata och
offentliga kapitalgivare är begränsad (se punkterna 107–116).
Rekommendation 5 – Skapa länkar till finansieringsinstrument
Kommissionen bör
regelbundet samla in information om det belopp och den typ av finansiering som
SMF-I-stödmottagarna behöver under genomförandet av innovationsprojektet,
öka medvetenheten bland stödmottagarna om att det finns olika
finansieringsinstrument på EU-nivå och nationell nivå, och ge råd om vilka av
dessa som skulle passa deras finansiella behov bäst,
identifiera och främja synergier med EU-stödda finansieringsinstrument för att
stödja SMF-I-stödmottagarna med deras anskaffande av kapital,
samarbeta med medlemsstaterna och nationella investeringsbanker för att främja
nationellt stödda finansieringsinstrument som kanske kan uppfylla de finansiella
behov som SMF-I-stödmottagarna har.
Måldatum för genomförande: 2022
Denna rapport antogs av revisionsrättens avdelning IV, med ledamoten
Alex Brenninkmeijer som ordförande, vid dess sammanträde i Luxemburg den
december 2019.
För revisionsrätten
Klaus-Heiner Lehne
ordförande
Bilagor
Bilaga I – Metod
Skrivbordsgranskning av offentliga dokument och kommissionens interna
dokument, såsom rättsliga grunder, riktlinjer, konsekvensbedömningar,
utvärderings- och övervakningsrapporter, förslag till rättsakter, meddelanden,
ståndpunktsdokument och andra relevanta handlingar.
Analytisk granskning av uppgifter från olika källor: CORDA, Business Objects,
resultattavlan för innovation och webbsökningar.
Onlineenkäter som skickades i mars 2019 till
—
—
—
stödmottagare och icke-utvalda sökande som fick en
spetskompetensstämpel, som valdes ut slumpmässigt, varav 71 % svarade
(88 % av de som fick stöd genom fas 2),
distansutvärderare som valdes ut slumpmässigt, med en svarsfrekvens
på 96 %,
nationella innovationsmyndigheter eller liknande organ, som alla svarade.
Informationsbesök till ministerier, innovationsmyndigheter, nationella
kontaktpunkter, EEN, stödmottagare och andra berörda intressenter i Bulgarien,
Danmark, Frankrike, Rumänien, Slovenien, Spanien och Förenade kungariket.
En panel med oberoende innovationsexperter inom olika områden.
Intervjuer med olika innovationsexperter med koppling till SMF-I, såsom
jurymedlemmar, medlemmar i den rådgivande gruppen av SMF-experter H2020
EAG och representanter för konsultföretag.
Deltagande i egenskap av observatörer i samband med jurypresentationer av
projekt (andra steget i urvalsprocessen till fas 2) och vid ett evenemang för
företagsaccelerationstjänster.
Intervjuer med kommissionspersonal vid GD Forskning och innovation,
GD Kommunikationsnät, innehåll och teknik, Easme och Genomförandeorganet
för forskning, liksom med EIB och EIF.
Bilaga II – Statistik
Finansiering per land (i milj. euro)
Spanien
Italien
Frankrike
Förenade kungariket
Tyskland
Sverige
Nederländerna
Danmark
Finland
Irland
Österrike
Belgien
Polen
Portugal
Ungern
Estland
Slovenien
Grekland
Tjeckien
Litauen
Kroatien
Slovakien
Malta
Lettland
Bulgarien
Cypern
Luxemburg
Rumänien
332,5
179,1
169,3
165,5
163,4
129,6
121,4
110,6
108,9
95,9
46,8
33,8
33,1
32,5
27,1
23,3
20,1
15,3
6,4
5,4
2,2
2,2
2,1
1,9
1,8
0,5
0,4
0,4
Finansiering per land,
i procent av den totala summan
Spanien
Italien
Frankrike
Förenade kungariket
Tyskland
Sverige
Nederländerna
Danmark
Finland
Irland
Österrike
Belgien
Polen
Portugal
Ungern
Estland
Slovenien
Grekland
Tjeckien
Litauen
Kroatien
Slovakien
Malta
Lettland
Bulgarien
Cypern
Luxemburg
Rumänien
2,6 %
1,8 %
1,8 %
1,8 %
1,5 %
1,3 %
1,1 %
0,8 %
0,3 %
0,3 %
0,1 %
0,1 %
0,1 %
0,1 %
0,1 %
0,0 %
0,0 %
0,0 %
0%
Förslag per land,
i procent av den totala summan
18,2 %
9,8 %
9,2 %
9,0 %
8,9 %
7,1 %
6,6 %
6,0 %
5,9 %
5,2 %
5%
%
%
Spanien
Italien
Frankrike
Förenade kungariket
Tyskland
Sverige
Nederländerna
Danmark
Finland
Irland
Österrike
Belgien
Polen
Portugal
Ungern
Estland
Slovenien
Grekland
Tjeckien
Litauen
Kroatien
Slovakien
Malta
Lettland
Bulgarien
Cypern
Luxemburg
Rumänien
Utvalda projekt per land,
i procent av den totala summan
Spanien
Italien
Frankrike
Förenade kungariket
Tyskland
Sverige
Nederländerna
Danmark
Finland
Irland
Österrike
Belgien
Polen
Portugal
Ungern
Estland
Slovenien
Grekland
Tjeckien
Litauen
Kroatien
Slovakien
Malta
Lettland
Bulgarien
Cypern
Luxemburg
Rumänien
7,1 %
9,9 %
7,6 %
5,6 %
4,9 %
4,7 %
3,6 %
3,0 %
2,8 %
1,8 %
1,9 %
2,7 %
1,9 %
1,4 %
1,4 %
0,7 %
0,5 %
0,7 %
0,2 %
0,5 %
0,1 %
0,3 %
0,3 %
0,2 %
0,2 %
0,2 %
0%
5%
%
8,9 %
6,7 %
4,3 %
4,3 %
3,0 %
3,5 %
2,1 %
1,7 %
1,7 %
3,3 %
2,4 %
3,3 %
1,4 %
2,0 %
1,6 %
1,1 %
0,7 %
0,6 %
1,1 %
0,1 %
0,9 %
1,8 %
0,4 %
0,2 %
0,9 %
5%
%
%
%
Framgångsgrad
per land
14,5 %
%
6,4 %
0%
%
17,8 %
17,9 %
%
21,4 %
Spanien
Italien
Frankrike
Förenade kungariket
Tyskland
Sverige
Nederländerna
Danmark
Finland
Irland
Österrike
Belgien
Polen
Portugal
Ungern
Estland
Slovenien
Grekland
Tjeckien
Litauen
Kroatien
Slovakien
Malta
Lettland
Bulgarien
Cypern
Luxemburg
Rumänien
%
Källa: Revisionsrätten på grundval av uppgifter från Easme.
5,6 %
7,6 %
7,6 %
7,8 %
8,9 %
7,9 %
10,6 %
7,0 %
9,6 %
11,6 %
7,0 %
4,0 %
8,0 %
4,0 %
4,8 %
3,1 %
3,5 %
2,0 %
3,0 %
4,3 %
2,3 %
1,2 %
4,3 %
1,2 %
0%
2%
4%
6%
8,3 %
7,1 %
7,3 %
6,6 %
% 10 % 12 % 14 %
Bilaga III – Europeiska innovationsrådet inom ramen för
Horisont Europa – från idé till förslag
—
I juni 2015, under ERA-konferensen ”A new start for Europe: Opening up to an
ERA of Innovation”, lanserade kommissionen idén om ett europeiskt
innovationsråd.
—
Kommissionen genomförde ett öppet samråd under våren 2016 för att bidra till
utformningen av pilotprojektet för ett europeiskt innovationsråd. Genom detta
offentliga samråd samlade kommissionen in intressenternas synpunkter om
disruptiv marknadsskapande innovation, om brister i det nuvarande landskapet
för innovationsstöd och om de potentiella befogenheterna för ett europeiskt
innovationsråd 39.
—
Den 13 juli 2016 anordnade kommissionen en workshop med över 100
intressenter från privat sektor, forskarvärlden och offentlig sektor för att
diskutera utfallet av det offentliga samrådet 40.
—
I november 2016 lanserade kommissionen initiativet för uppstartsföretag och
expanderande företag, som syftar till att sammanföra en mängd befintliga och
nya åtgärder under samma paraply för att stödja uppstartsföretag och företag
som vill skala upp sin verksamhet 41.
Ideas for an EIC, sammanfattning av svaren på förfrågan om idéer, 2016.
Ideas for an EIC – sammanfattning av en valideringsworkshop med intressenter som
anordnades den 13 juli 2016.
COM(2016) 733 final, meddelande, Europas nästa ledare – initiativet för uppstartsföretag
och expanderande företag, november 2016.
—
Kommissionen inrättade EIC:s högnivågrupp av innovatörer (EIC High Level Group
of Innovators) i januari 2017, som fick i uppdrag att tillhandahålla stöd till
utvecklingen av Europeiska innovationsrådet. Denna grupp, som bestod av
företagare, investerare och innovationsexperter, möttes sex gånger mellan
mars 2017 och december 2018 och tog fram en komplett uppsättning
rekommendationer i januari 2018 42.
—
Den 7 juni 2018 lade kommissionen fram ett förslag till Europaparlamentets och
rådets förordning om inrättande av Horisont Europa. 43 En konsekvensbedömning
åtföljde förslaget 44.
Europe is back: Accelerating breakthrough innovation, EIC:s högnivågrupp, januari 2018.
COM(2018) 435 final, Förslag till förordning om inrättande av Horisont Europa, juni 2018.
SWD(2018) 307 final, arbetsdokument från kommissionens avdelningar,
konsekvensbedömning, juni 2018.
Akronymer och förkortningar
BNP: bruttonationalprodukt.
EAG: den rådgivande gruppen av SMF-experter.
Easme: Genomförandeorganet för små och medelstora företag.
EEN: Enterprise Europe Network.
EIB: Europeiska investeringsbanken.
EIC: Europeiska innovationsrådet.
EIF: Europeiska investeringsfonden.
FoU: forskning och utveckling.
GD Forskning och innovation: kommissionens generaldirektorat för forskning och
innovation.
H2020: Horisont 2020.
it: informationsteknik.
SBIR: programmet för innovation och forskning i små företag (USA).
SMF: små och medelstora företag.
SMF-I: EU:s instrument för små och medelstora företag.
Ordlista
associerat land: ett tredjeland som är part i ett internationellt avtal med Europeiska
unionen; associerade länder till ramprogrammet Horisont 2020 deltar på samma villkor
som juridiska enheter från EU:s medlemsstater.
banbrytande innovation: en produkt, tjänst eller process som introducerar en ny
teknik eller en ny affärsmodell som leder till ett paradigmskifte och innebär betydande
konkurrensfördelar.
blandad finansiering: en kombination av bidrag och lån eller kapital från offentliga
eller privata källor.
deltagarportal: den enda onlineportalen för sökande och stödmottagare inom ramen
för Horisont 2020 för att identifiera finansieringsmöjligheter, få tag på dokument och
få vägledning, lämna in förslag och för papperslös hantering av bidrag och expertavtal;
se http://ec.europa.eu/research/participants/portal.
disruptiv innovation: en produkt, tjänst eller process som splittrar de befintliga
marknaderna genom att tränga undan ledande företag och tekniker och tillämpa nya
värderingar.
europeisk resultattavla för innovation: en jämförande analys av hur EUmedlemsstaterna, andra europeiska länder och regionala grannar presterar när det
gäller innovation.
finansieringsinstrument: ekonomiskt stöd från EU-budgeten i form av investeringar av
eget kapital, investeringar av kapital likställt med eget kapital, lån eller garantier eller
andra riskdelningsinstrument.
förslagsinfordran: ett dokument som efterlyser ansökningar från potentiella
stödmottagare, som offentliggörs av en offentlig enhet som tillkännager sin avsikt att
finansiera projekt som uppfyller angivna syften.
inlämningsdatum: det datum som förslagen senast måste lämnas in för en särskild
finansieringsomgång.
nationell kontaktpunkt: en nationell enhet som inrättats och finansieras av
regeringarna i EU:s medlemsstater eller stater som är associerade till ett ramprogram
för forskning för att tillhandahålla stöd på plats och vägledning till de som ansöker om
och får stöd från Horisont 2020.
stödmottagare: en fysisk eller juridisk person som får ett bidrag eller lån från EU:s
budget.
KOMMISSIONENS SVAR PÅ EUROPEISKA REVISIONSRÄTTENS SÄRSKILDA
RAPPORT
SMF-INSTRUMENTET I PRAKTIKEN: ETT ÄNDAMÅLSENLIGT OCH INNOVATIVT
PROGRAM SOM STÅR INFÖR UTMANINGAR”
I. Instrumentet för små och medelstora företag (nedan kallat SMF-instrumentet) är den första
stödordningen någonsin inom ramprogrammet för forskning som är inriktad på innovativa små och
medelstora företag och som genomförs via ett genomförandeorgan. Små och medelstora företag vars
stöd släpat efter i tidigare ramprogram har i stor utsträckning anslutit sig till detta nya stödsystem
som, med tiden, har finjusterats för att bättre motsvara deras faktiska behov. Framgången med den
första omgången av Europeiska innovationsrådets (nedan kallat EIC) pilotprogram Accelerator visar
att den väg som kommissionen slagit in på ligger i linje med förväntningarna hos innovativa små och
medelstora företag.
INLEDNING
Kommissionen har genomfört tester av ekonomiskt stöd till projekt genom finansiering med eget
kapital från och med oktober 2019.
IAKTTAGELSER
Medlemmar i kommittén för tillgång till riskfinansiering och programkommittén för små och
medelstora företag, som ofta också är nationella kontaktpunkter, har regelbundet informerats om de
ändringar som införts i SMF-instrumentet.
Dessutom gjordes informationskampanjer om sådana förändringar av GD Forskning och innovation
och genomförandeorganet för små och medelstora företag (nedan kallat Easme) för att öka
medvetenheten hos de berörda parterna, inklusive de nationella kontaktpunkterna och Enterprise
Europe Network (EEN).
SMF-instrumentet är inriktat på alla typer av innovativa små och medelstora företag som visar en
stark strävan att utvecklas, växa och internationaliseras.
I linje med den nya kommissionsordförandens politiska prioriteringar planerar man att genomföra en
särskild ansökningsomgång för EIC:s Accelerator-program för 2020, med förbehåll för godkännande
från kommittén för det strategiska programmet.
Kommissionen påpekar att denna risk har tagits upp i EIC-pilotprojektet från och med 2019.
Dessutom betonas att det finns en stor klyfta mellan uppfattningen hos stödmottagare inom ramen för
SMF-I och den verkliga situationen när det gäller att skaffa fram pengar från riskkapital eller
affärsänglar, där det visar sig att framgången är tämligen begränsad.
Kommissionen understryker att den har gjort stora ansträngningar för att främja EIC:s (förstärkta)
pilotprogram och anordna seminarier för SMF-I vid olika teknikkonferenser runtom i Europa (bl.a.
Slush, Wolves Summit, Smart City). De ändringar som infördes genom det förbättrade EICpilotprojektet kommunicerades via kampanjturnéer och särskilda evenemang som anordnats i alla
medlemsstater.
Sedan Horisont 2020 inleddes har mer än 65 uppsökande evenemang anordnats i medlemsstater och
associerade länder. Kommissionens informationskampanj i medlemsstaterna, som anordnades i
samarbete med de nationella kontaktpunkterna, intensifierades under 2019 med deltagandet av små
och medelstora företag. Kommissionen inledde därefter en omgång nationella och regionala samråd
med berörda parter, som pågår i medlemsstaterna sedan juni 2019, för att gemensamt utforma
genomförandet av Horisont Europa, där nästa strategi för små och medelstora företag kommer att
fastställas.
Kommissionen anser att samordnings- och stödinsatsen Access4SME har bidragit till att öka
medvetenheten bland de nationella kontaktpunkterna och EEN i anslutning till att förändringar har
gjorts i utformningen av SMF-instrumentet.
Easme behövde faktiskt förnya 25 % av gruppen av utvärderare på årsbasis för att följa H2020reglerna.
Som svar på behovet av utbildning av nytillkomna har Easme sedan 2018 arrangerat expertdagar i
Bryssel och bjudit in både erfarna och nya experter till att delta i fortbildning och skapa synergier.
På grundval av synpunkterna från jurymedlemmarna införde kommissionen i oktober 2019 en
praxis som innebär att jurymedlemmarna har två veckor på sig att grundligt gå igenom förslagen.
För att komma till rätta med det problem som revisionsrätten påpekar i denna punkt har
kommissionen infört ett förfarande för tillbörlig aktsamhet i EIC:s förstärkta pilotprojekt. Inom ramen
för det förstärkta EIC-pilotprojektet som erbjuder blandad finansiering har man från och med oktober
begärt mer ingående information från de sökande med avseende på ägande, immateriella
rättigheter och gruppsammansättning. Dessa aspekter bedöms nu av utvärderarna via kontakter på
distans och genom intervjuer.
Även om det inte föreskrivs i den rättsliga grunden för SMF-instrumentet och med förbehåll för
godkännande av den berörda programkommittén, kan kommissionen komma att föreslå ett förfarande
som begränsar antalet förnyade inlämningar.
Kommissionen betonar att starten av företagsaccelerationstjänsterna föregicks av grundliga
förberedelser och ett öppet upphandlingsförfarande.
Easme samlar in information om ytterligare finansieringsbehov hos vissa stödmottagare, under
och efter genomförandeperioden för bidraget, något som görs genom flera kanaler (ansökningar till
BAS-investerarevenemang och företagsprofil i Scaleup-verktyget för matchning mellan investerare).
Från och med inlämningsfristen oktober 2019 måste företagen dessutom ange hur de avser att
finansiera all nödvändig utvecklingsverksamhet till dess att marknadsinträde sker, utöver det begärda
bidraget och/eller eget kapital. Detta inbegriper uppgifter om både de belopp som krävs och källor till
potentiell finansiering.
Kommissionen har börjat ta itu med den fråga som revisionsrätten nämner i denna punkt genom
genomförandet av EIC:s förstärkta pilotprojekt 2019.
SLUTSATSER OCH REKOMMENDATIONER
Att nå ut till och kommunicera med berörda parter är en av kommissionens huvudprioriteringar
för ett sunt genomförande av de nuvarande och framtida ramprogrammen. Kontaktskapande
verksamhet avseende formerna för genomförandet av Horisont 2020 anordnas regelbundet i
medlemsstater och associerade länder. Ytterligare en rad evenemang i medlemsstaterna är inriktade på
Horisont Europa.
Rekommendation 1 – Förbättra kommunikationsstrategin och stödet till de nationella
kontaktpunkterna, i synnerhet för de medlemsstater som har lägst deltagande
Kommissionen godtar rekommendationen.
Kommissionen avser att planera en ny strategi i enlighet med rekommendationen från januari
för Horisont Europa.
Rekommendation 2 – Förbättra urvalsförfarandet
Kommissionen godtar rekommendationen.
Kommissionen har genomfört denna rekommendation från och med den utvärdering som inleddes i
oktober 2019 genom att skicka förslagen två veckor i förväg. Från och med mars 2020 kommer
dessutom de externa experterna att ha 0,5 dagar på sig att utvärdera ett förslag, jämfört med 0,3 dagar
till och med januari 2020.
Kommissionen avser att genomföra en ny strategi i enlighet med rekommendationen från januari
Kommissionen anger att den redan offentliggör framgångsgraden per inlämnat förslag och
samtycker till att även lägga till framgångsgraden per projektförslag.
Rekommendation 3 – Ersätt fas 1 och bygg vidare på fas 2-stödet till små och medelstora
företag
Kommissionen godtar rekommendationen.
En del medlemsstater under ledning av Tjeckien har inrättat en informell arbetsgrupp för att kopiera
fas 1, som finansieras på nationell nivå men fortfarande omfattas av en central EU-utvärdering.
Kommissionen kan komma att föreslå att de ska stödjas i sitt samordningsarbete genom ett särskilt
bidrag.
I det partiella allmänna avtalet om Horisont Europa förutses en fortsättning av systemet med enbart
bidrag inom EIC:s Accelerator, med en budget motsvarande den för Horisont 2020, samtidigt som
budgeten för EIC:s Accelerator främst bör användas för blandfinansiering.
Rekommendation 4 – Förbättra företagsaccelerationstjänsterna
Kommissionen godtar rekommendationen, inom ramen för de resurser som är tillgängliga för
efterföljaren till SMF-instrumentet inom ramen för nästa fleråriga budgetram.
När det gäller att öka stödmottagarnas medvetenhet har EIB och EIF genomfört en bred
informationskampanj med avseende på InnovFin-finansieringsinstrumenten i alla medlemsstater
mellan 2014 och 2016, och därvid utvecklat kontakter med många små och medelstora företag, trots
att kampanjen inte riktade sig specifikt till företag som mottar stöd genom SMF-instrumentet. En
informationskampanj om EIC:s förstärkta pilotprogram som lanserades under våren 2019 ökade
medvetenheten hos potentiella stödmottagare om möjlig finansiering med eget kapital genom EIC:s
Accelerator.
Kommissionen har också börjat samla in uppgifter från ansökningsprocessen från inlämningsfristen
oktober 2019 om de finansiella behoven, inbegripet bidrag och eget kapital hos företag som ansöker
för att ha möjlighet att framgångsrikt expandera.
Rekommendation 5 – Skapa länkar till finansiella instrument
Kommissionen godtar rekommendationen.
Bidrags- och investeringsavtalen kommer att regelbundet övervaka de finansiella behoven under hela
projektets genomförande och under expansionsfasen.
Kommissionen godtar rekommendationen.
Kommissionen kommer att fortsätta sin informationsverksamhet.
Kommissionen godtar rekommendationen.
I det partiella allmänna avtalet om Horisont Europa förutses möjligheten för stödmottagare att ansöka
om eget kapital först från och med 2021.
Kommissionen godtar delvis rekommendationen.
Med hänsyn till att rekommendationen även berör medlemsstater, kan kommissionen endast åta sig att
följa den efter bästa förmåga.
Kommissionen kommer att bidra till att öka medlemsstaternas och nationella utvecklingsinstitutioners
medvetenhet genom den berörda programkommittén.
Införandet av spetskompetensstämpeln för framgångsrika förslag som inte kunde beviljas bidrag ur
SMF-instrumentet var ett första försök att skapa synergier med nationella ekosystem som stöder
innovation.
Granskningsteam
I våra särskilda rapporter redovisar vi resultatet av våra revisioner av EU:s politik och
program eller av förvaltningsteman kopplade till specifika budgetområden. För att
uppnå så stor effekt som möjligt väljer vi ut och utformar granskningsuppgifterna med
hänsyn till riskerna när det gäller prestation eller regelefterlevnad, storleken på de
aktuella intäkterna eller kostnaderna, framtida utveckling och politiskt intresse och
allmänintresse.
Denna effektivitetsrevision utfördes av revisionsrättens avdelning IV
marknadsreglering och en konkurrenskraftig ekonomi, där ledamoten
Alex Brenninkmeijer är ordförande. Han ledde revisionsarbetet med stöd av
Raphael Debets (kanslichef), John Sweeney (förstechef), Juan Antonio Vazquez Rivera
(uppgiftsansvarig) och Alvaro Garrido-Lestache Angulo, Wayne Codd och
Marco Montorio (revisorer).
Från vänster till höger: John Sweeney, Marco Montorio, Raphael Debets, Juan Antonio
Vazquez Rivera, Wayne Codd , Alex Brenninkmeijer, Alvaro Garrido-Lestache Angulo.
Tidslinje
Händelse
Datum
Revisionsplanen antogs/Revisionen inleddes
2019
Den preliminära rapporten skickades till kommissionen
(eller andra revisionsobjekt)
2019
Den slutliga rapporten antogs efter det kontradiktoriska
förfarandet
2019
Svaren från kommissionen (eller från ett annat revisionsobjekt)
hade tagits emot på alla språk
2020
UPPHOVSRÄTT
© Europeiska unionen 2020.
Europeiska revisionsrättens policy för vidareutnyttjande av handlingar tillämpas genom Europeiska
revisionsrättens beslut nr 6-2019 om öppen datapolitik och vidareutnyttjande av handlingar.
Om inget annat anges (t.ex. i enskilda meddelanden om upphovsrätt) omfattas revisionsrättens
innehåll som ägs av EU av den internationella licensen Creative Commons Erkännande 4.0 (CC BY 4.0).
Det innebär att vidareutnyttjande är tillåtet under förutsättning att ursprunget anges korrekt och att
det framgår om ändringar har gjorts. Vidareutnyttjas materialet får handlingarnas ursprungliga
betydelse eller budskap inte förvanskas. Revisionsrätten bär inte ansvaret för eventuella konsekvenser
av vidareutnyttjande.
När enskilda privatpersoner kan identifieras i ett specifikt sammanhang, exempelvis på bilder av
revisionsrättens personal, eller om arbete av tredje part används, måste tillstånd inhämtas med
avseende på de ytterligare rättigheterna. Om tillstånd beviljas upphävs det allmänna godkännande
som nämns ovan och eventuella begränsningar av materialets användning måste tydligt anges.
För användning eller återgivning av innehåll som inte ägs av EU kan tillstånd behöva inhämtas direkt
från upphovsrättsinnehavarna. Programvara eller handlingar som omfattas av immateriella rättigheter,
till exempel patent, varumärkesskydd, mönsterskydd samt upphovsrätt till logotyper eller namn,
omfattas inte av revisionsrättens policy för vidareutnyttjande eller av licensen.
EU-institutionernas webbplatser inom domänen europa.eu innehåller länkar till webbplatser utanför
den domänen. Eftersom revisionsrätten inte kontrollerar dem uppmanas du att ta reda på vilken
integritetspolicy de tillämpar.
Användning av Europeiska revisionsrättens logotyp
Användningen av Europeiska revisionsrättens logotyp måste först godkännas av Europeiska
revisionsrätten.
PDF
HTML
ISBN: 978-92-847-4153-3
ISBN: 978-92-847-4133-5
ISSN: 1977-5830
ISSN: 1977-5830
doi: 10.2865/841285
doi: 10.2865/1789
QJ-AB-19-025-SV-N
QJ-AB-19-025-SV-Q
Med 3 miljarder euro i anslag för 2014–2020 ska EU:s SMFinstrument stödja innovation i små och medelstora företag och
uppstartsföretag genom att avhjälpa bristen på finansiering och
öka kommersialiseringen av forskningsresultat.
Vi bedömde om SMF-instrumentet leder till de förväntade
fördelarna. Vi drog den övergripande slutsatsen att instrumentet
ger ändamålsenligt stöd till små och medelstora företag när de
utvecklar sina innovationsprojekt. EU:s varumärke hjälper
dessutom företagen att locka till sig ytterligare investeringar.
Kommissionen förvaltar instrumentet på ett kompetent sätt. Vi
rekommenderar dock förbättringar när det gäller inriktningen på
stödmottagare, geografisk spridning och urval av projekt. Mer kan
också göras för att attrahera ytterligare finansiering som skulle
hjälpa till att lansera innovationsprojekt på marknaden.
SMF-instrumentet har omformats inför perioden 2021–2027 som
en del av Europeiska innovationsrådet (EIC), och våra
rekommendationer gäller framför allt aspekter av utformningen
som bör bevaras, förbättringar i urvalet av projekt, utökade
företagsaccelerationstjänster och skapandet av synergier med
andra finansieringsinstrument.
Revisionsrättens särskilda rapport i enlighet med artikel 287.4
andra stycket i EUF-fördraget.
Särskild rapport
EU:s investeringar i kulturplatser:
ökat fokus och bättre samordning
behövs
Innehållsförteckning
Punkt
Sammanfattning
I–VIII
Inledning
01–11
Revisionens inriktning och omfattning samt
revisionsmetod
12–16
Iakttagelser
17–93
Den befintliga ramen för EU:s investeringar i kulturplatser saknar
fokus, och samordningen är begränsad
17–51
Den strategiska ramen för EU:s insatser för kultur är komplex och
återspeglas endast delvis i EU:s finansiering
17–24
Kommissionen har utvecklat flera initiativ som kan främja kulturplatser,
men samordningen med finansieringsarrangemang är begränsad
25–36
Eruf är ett instrument för att strukturera medlemsstaternas investeringar i
kulturplatser, men sådana investeringar behandlas inte som en prioritering
för Eruf
37–51
Varierande ändamålsenlighet och hållbarhet hos de granskade
Eruf-projekten
52–93
De slutförda, granskade projekten var operativa, deras mål var för det mesta
ekonomiska och det gick inte alltid att säga om de hade uppnåtts
55–67
Otillräcklig uppmärksamhet ägnas åt kulturplatsers hållbarhet
68–93
Slutsatser och rekommendationer
94–105
Bilagor
Bilaga I – Översikt över offentliga utgifter för kulturella tjänster
Bilaga II – Översikt över EU-fonder med kulturella mål
Bilaga III – Lista över granskade insatsområden och tillhörande
operativa program
Bilaga IV – Lista över granskade projekt
Bilaga V – Översikt över de 21 granskade urvalsförfarandena
Bilaga VI – Lista över de viktigaste policydokumenten avseende
kulturplatser
Bilaga VII – Viktigaste kännetecken för europeiska
kulturarvsmärket, världsarvslistan och kulturvägar
Bilaga VIII – Utveckling av Eruf-ramen för investeringar i
kulturplatser
Bilaga IX – Viktigaste målen för insatsområdena i urvalet och
mätning av dem med resultatindikatorer
Akronymer och förkortningar
Ordlista
Kommissionens svar
Granskningsteam
Tidslinje
Sammanfattning
I De flesta européer anser att kulturarvet är viktigt för dem personligen liksom för
deras kommun, region och land samt för EU i stort. Kultur är ett vitt begrepp som
inbegriper olika aktiviteter. I den här särskilda rapporten avses med ”kulturplatser”
den fysiska infrastruktur där européer kan uppleva kultur.
II EU:s kulturella ram definieras primärt i fördragen. Där anges som överordnat mål
att EU ska respektera rikedomen hos sin kulturella mångfald och sörja för att det
europeiska kulturarvet skyddas och utvecklas. Kultur är huvudsakligen
medlemsstaternas behörighet. Unionen kan endast uppmuntra till samarbete mellan
medlemsstater och stödja eller komplettera deras insatser.
III Vi bedömde ändamålsenligheten och hållbarheten i Eruf-investeringar i
kulturplatser genom att bedöma hur lämplig EU:s kulturella ram är, hur den samordnas
med finansieringsarrangemang och hur Eruf-finansieringen genomförs.
IV Revisionen var inriktad på de ekonomiska, sociala och kulturella effekterna av
investeringarna och på kulturplatsernas finansiella och fysiska hållbarhet. Vi granskade
kommissionens arbete och bedömde 27 projekt i sju medlemsstater. Vi intervjuade
även experter på området.
V Den samlade slutsatsen av revisionen är att den nuvarande ramen saknar fokus och
behöver samordnas bättre för att säkerställa att Eruf-investeringarna i kulturplatser
blir ändamålsenliga och hållbara. Vi gjorde nedanstående iakttagelser.
VI Vad beträffar ramen för EU:s investeringar i kulturplatser:
o
Kultur behandlas inte i kommissionens övergripande Europa 2020-strategi. EU:s
grundläggande strategiska ram för kultur är komplex och återspeglas endast
delvis i EU:s finansiering. Enligt kommissionen är det fortfarande en utmaning att
omvandla EU-målen till politiska beslut på medlemsstatsnivå.
o
Kommissionen har utvecklat flera initiativ som kan främja kulturplatser, men EU:s
kulturinitiativ har begränsad effekt på stödmottagares tillgång till EU-medel. Erufförordningen innehåller inga bestämmelser som gagnar kulturplatser som deltar i
EU:s kulturinitiativ. Samordningen mellan EU:s fonder när det gäller investeringar
i kulturplatser är också begränsad.
o
På EU-nivå finansieras infrastrukturinvesteringar framför allt genom Eruf, som för
omkring en tredjedel av medlemsstaterna är en viktig källa till finansiering av
offentliga investeringar i kulturplatser. Men Eruf prioriterar inte investeringar i
kulturplatser utan stöder ett annat fördragsmål: främjandet av social och
ekonomisk sammanhållning. På nationell nivå fann vi exempel på
medlemsstatsinitiativ som gick ut på att finansiera kulturplatser med privata
medel.
VII Vad beträffar ändamålsenligheten och hållbarheten hos de granskade Eruf-
projekten:
o
Trots EU:s ambition att öka kulturinsatsernas sociala effekter är målen för Erufs
operativa program och projekt mestadels ekonomiska. I de operativa program
som vi granskade ägnades minst uppmärksamhet åt kulturella aspekter, och de
flesta förvaltande myndigheter betraktar inte ens kulturella aspekter som ett
kriterium när de väljer ut projekt.
o
Projektens prestation kunde endast bedömas för vissa av de slutförda, granskade
projekten. Projekten var operativa, men vi fann flera brister i urvalet och
rapporteringen av indikatorer, vilket begränsar möjligheten att använda de
rapporterade uppgifterna för att dra slutsatser om projektens prestation.
o
Varken Eruf eller Kreativa Europa kan finansiera bevarandet av utsatta
kulturplatser om inte arbetet har direkta ekonomiska och sociala effekter.
Skapandet av ekonomiska effekter, ofta genom strategier för turismfrämjande,
kan vara kontraproduktivt för bevarandet av kulturarvsplatser.
o
De granskade kulturplatserna är i allmänhet beroende av offentliga subventioner
för sin drift och finansiering av investeringskostnader. Den nuvarande
finansieringsramen ger inte tillräckliga incitament till inkomstgenerering. Erufkraven på inkomstgenererande projekt innebär att ju högre nettoinkomster som
projektet genererar, desto mindre blir EU-stödet. De urvalsförfaranden som vi
granskade gav sällan incitament till inkomstgenererande verksamhet.
VIII För att säkerställa sund ekonomisk förvaltning i samband med investeringar i
kulturplatser rekommenderar vi att kommissionen
förbättrar den nuvarande strategiska ramen för kultur i enlighet med de
befogenheter som anges i fördragen,
uppmuntrar användning av privata medel för att skydda Europas kulturarv,
stärker den finansiella hållbarheten för kulturplatser som finansieras av Eruf,
vidtar mer specifika åtgärder för att bevara kulturarvsplatser.
Inledning
Kultur och kulturplatser
De flesta européer anser att kulturarvet är viktigt för dem personligen liksom för
deras kommun, region och land samt för EU i stort 1. Kultur är också en resurs.
Kommissionen har identifierat kultur som en drivkraft för tillväxt och jobb,
möjliggörare av social integration och en tillgång för att stärka EU:s internationella
relationer 2. Enligt statistik från Eurostat sysselsatte kultursektorn 8,7 miljoner
människor i EU 2018 eller 3,8 % av den totala arbetskraften 3.
Kultur är ett vitt begrepp som inbegriper olika aktiviteter (t.ex. hantverk, konst
och audiovisuell verksamhet) inom olika ekonomiska sektorer (t.ex. tillverkning,
tjänster och kommunikation). I den här särskilda rapporten avses med ”kulturplatser”
den fysiska infrastruktur där européer kan uppleva kultur. Vi skiljer mellan
kulturarvsplatser (gamla historiska platser) och ny kulturell infrastruktur (nya
byggnader som används för att främja konst, musik, teater etc.).
Beslutsfattandet på EU-nivå tog fart 2017 när EU:s ledare uppmanades att göra
mer inom områdena utbildning och kultur 4. På senare tid har Europeiska rådet i sin nya
strategiska agenda för 2019–2024 åtagit sig att ”investera i kultur och i vårt kulturarv,
vilka är centrala för den europeiska identiteten” 5.
Politisk ram
I fördragen anges att EU ”ska respektera rikedomen hos sin kulturella
mångfald och sörja för att det europeiska kulturarvet skyddas och utvecklas” 6, och att
EU ska stödja kultur i medlemsstaterna 7. Fördragen anger också på vilka områden EU
ska vidta åtgärder (spridning av kulturen, kulturarv, icke-kommersiellt kulturutbyte,
Cultural Heritage, särskild Eurobarometer, nr 466, enkät gjord på begäran av Europeiska
kommissionen, december 2017.
Meddelande från kommissionen om en europeisk agenda för en kultur i en alltmer
globaliserad värld, KOM(2007) 242 slutlig, 10.5.2007.
Eurostat, Culture statistics, fjärde upplagan, 2019, s. 64.
Europeiska rådets möte, 14 december 2017, EUCO 19/1/17.
En ny strategisk agenda 2019–2024, Europeiska rådet.
Artikel 3.3 i EU-fördraget.
Artikel 167.1 i EUF-fördraget.
konstnärligt och litterärt skapande och externt samarbete). De fastställer också ett
allmänt krav på insatser på andra politikområden för att beakta kulturella aspekter,
vilket kallas ”integrering” 8.
EU har ingen lagstiftningsbehörighet på kulturområdet. Ansvaret för
beslutsfattandet på detta område ligger hos medlemsstaterna. År 2017 anslog
medlemsstaterna 1 % av sina offentliga utgifter till kulturella tjänster, vilket innebär att
euro per EU-medborgare gick till stöd för kulturella aktiviteter. Av det beloppet
användes omkring 15 % till kulturella investeringar (dvs. förvärv, skapande eller
restaurering av kulturtillgångar, inbegripet fysiskt arbete på kulturplatser). Bilaga I
innehåller närmare uppgifter om de offentliga utgifterna för kulturella tjänster och
kulturella investeringar i EU.
Ramen för EU-samarbete på kulturområdet fastställs av kommissionen i den
europeiska agendan för kultur. Den första agendan antogs 2007 9. År 2018 antog
kommissionen en ”ny agenda för kultur” 10. Den nya agendan har följande tre
strategiska mål:
—
Den sociala dimensionen – att ta tillvara den inneboende styrkan hos kultur och
kulturell mångfald för att främja social sammanhållning och välfärd genom att
uppmuntra till kulturellt deltagande, rörlighet bland konstnärer och skydd av
kulturarv.
—
Den ekonomiska dimensionen – att stödja sysselsättning och tillväxt i de kulturella
och kreativa sektorerna genom att främja konst och kultur inom utbildning,
främja relevant kompetens och uppmuntra innovation inom kulturen.
—
Den externa dimensionen – att stärka de internationella kulturella förbindelserna
genom att till fullo utnyttja kulturens potential att gynna hållbar utveckling och
fred.
Den nya agendan fastställer åtgärder som kommissionen ska vidta och uppmanar
medlemsstaterna att ta upp vissa frågor. Medlemsstaterna anger sina prioriteringar för
Artikel 167.4 i EUF-fördraget: ”Unionen ska beakta de kulturella aspekterna då den handlar
enligt andra bestämmelser i fördragen, särskilt för att respektera och främja sin kulturella
mångfald”.
Meddelande från kommissionen om en europeisk agenda för en kultur i en alltmer
globaliserad värld, KOM(2007) 242 slutlig, 10.5.2007.
Kommissionens meddelande En ny europeisk agenda för kultur, COM(2018) 267 final,
2018.
EU-samarbetet om kultur och arbetsmetoder genom arbetsplaner för kultur som antas
av ministerrådet. Den senaste arbetsplanen omfattar perioden 2019–2022 11.
Hållbarhet och kultur
EU och medlemsstaterna deltar också aktivt i multilaterala forum och
organisationer som arbetar med kultur- och kulturarvspolitik, till exempel Europarådet
och Unesco. Nu senast åtog sig EU:s medlemsstater att försöka uppnå de mål för
hållbar utveckling som tagits fram av Unesco 12 och på så vis förstärka det mål för
hållbar utveckling som fastställs i fördragen 13. Rådet har också identifierat kulturarvets
hållbarhet som en prioritering i den nuvarande arbetsplanen för kultur 2019–2022.
Styrning vid kommissionen
För närvarande ansvarar kommissionens generaldirektorat för utbildning,
ungdom, idrott och kultur (GD Utbildning, ungdom, idrott och kultur) för att utarbeta
och genomföra kulturrelaterad politik. Till stöd för EU:s kulturpolitiska beslutsfattande
förvaltar kommissionen programmet Kreativa Europa, som är den enda fonden som
uteslutande är inriktad på EU:s kulturella och kreativa näringar 14.
Kulturrelaterade infrastrukturinvesteringar kan endast EU-finansieras inom
ramen för de europeiska struktur- och investeringsfonderna (ESI-fonderna). Bland ESIfonderna är Eruf 15 den främsta källan till EU-finansiering av investeringar i
kulturplatser. Eruf genomförs av kommissionen och medlemsstaterna genom delad
förvaltning. Det betyder att partnerskapsöverenskommelserna och de operativa
programmen inom Eruf utarbetas av medlemsstaterna och måste godkännas av
kommissionen.
Rådets slutsatser om arbetsplanen för kultur 2019–2022 (EUT C 460, 21.12.2018, s. 12).
Att förändra vår värld: Agenda 2030 för hållbar utveckling, antagen av FN den
september 2015.
Artikel 3.3 i EU-fördraget.
Europaparlamentets och rådets förordning (EU) nr 1295/2013 av den 11 december 2013
om inrättande av programmet Kreativa Europa (2014–2020), EUT L 347, 20.12.2013, s. 221.
Kreativa Europa omfattar även den audiovisuella sektorn.
Europaparlamentets och rådets förordning (EU) nr 1301/2013 av den 17 december 2013
om Europeiska regionala utvecklingsfonden och om särskilda bestämmelser för målet
Investering för tillväxt och sysselsättning (EUT L 347, 20.12.2013, s. 289).
Till följd av principen om integrering är även andra EU-fonder tillgängliga för
kulturrelaterade projekt både inom och utanför EU. Det innebär att flera
generaldirektorat också är inblandade i det faktiska genomförandet av den kulturella
strategiramen via annan EU-politik och andra finansieringsinstrument (se bilaga II).
Revisionens inriktning och omfattning
samt revisionsmetod
Med tanke på den ökade uppmärksamhet som kultur röner på EU-nivå beslutade
vi att utföra en revision av hållbarheten och ändamålsenligheten i EU:s investeringar i
kulturplatser, det vill säga förvärv, återställande och skapande av ny kulturell
infrastruktur och kulturarvsplatser. Därför granskade vi den viktigaste EU-fond som
finns tillgänglig för sådana investeringar (Eruf) och bedömde nedanstående aspekter.
Del 1: Lämplighet hos EU:s kulturella ram och samordning med
finansieringsarrangemang för investeringar i kulturplatser
—
Lämpligheten hos den strategiska och rättsliga ram som har införts på EU-nivå för
EU-finansierade investeringar i kulturplatser.
—
Samordningen mellan de finansiella och politiska instrumenten i kommissionens
initiativ, särskilt med Kreativa Europa och Ejflu.
—
Samordningen av Eruf-finansiering med andra EU-fonder.
Del 2: Genomförande av Eruf-finansiering
—
Det stöd och den vägledning som kommissionen ger medlemsstaterna när de
antar partnerskapsöverenskommelser och operativa program för att säkerställa
att finansieringen av kulturplatser leder till ändamålsenliga och hållbara resultat.
—
Ändamålsenligheten och hållbarheten i resultaten av Eruf-projekt om
kulturplatser.
Revisionen var inriktad på de ekonomiska, sociala och kulturella effekterna av
Eruf-investeringar i kulturplatser och på platsernas hållbarhet i ekonomiskt och fysiskt
hänseende. Den omfattade programperioderna 2007–2013 och 2014–2020 inom
målet Investering för tillväxt och sysselsättning samt förslaget till utformning av
programperioden efter 2020.
På EU-nivå granskade vi det arbete som generaldirektoratet med ansvar för kultur
(GD Utbildning, ungdom, idrott och kultur) och generaldirektoratet med ansvar för Eruf
(GD Regional- och stadspolitik) hade utfört. På medlemsstatsnivå gjorde vi följande:
o
Vi besökte tre medlemsstater (Italien, Polen och Portugal) och utförde
skrivbordsgranskningar av mer begränsad omfattning för ytterligare fyra
medlemsstater (Kroatien, Frankrike, Tyskland och Rumänien). Vi valde dessa
medlemsstater eftersom de är bland de största mottagarna av Eruf-stöd för
investeringar i kulturplatser.
o
Vi bedömde 14 operativa program (i bilaga III finns en lista över de granskade
operativa programmen).
o
Vi granskade 27 projekt, varav 15 på plats och 12 genom skrivbordsgranskningar
(se tabell 1 och bilaga IV). Projekten valdes ut utifrån en rad olika kriterier:
belopp som använts eller anslagits, typ av plats (kulturarvsplats eller ny kulturell
infrastruktur), förekomst av utmärkelser och deltagande i EU-initiativ. Vi
genomförde även en enkät bland stödmottagarna i alla dessa projekt som
samtliga stödmottagare besvarade. Vi granskade även 21 urvalsförfaranden
(se bilaga V).
Tabell 1 – Antal och typer av projekt som ingick i revisionen
2007–2013
Kulturarvsplatser
Antal projekt
2014–2020
Ny kulturell infrastruktur
Totalt
Kulturarvsplatser
Projekt som besöktes på plats i
-
Italien
-
Polen
-
Portugal
Granskade projekt som gällde
-
Tyskland
e.t.
-
Frankrike
e.t.
-
Kroatien
e.t.
-
Rumänien
e.t.
Källa: Revisionsrätten.
Slutligen intervjuade vi tjänstemän vid internationella organisationer (Unescos
världsarvscentrum, Europarådets kulturvägar och ICOMOS) och den icke-statliga
organisationen Europa Nostra samt 11 nationella experter i de tre besökta
medlemsstaterna för att få en bättre bild av de behov och utmaningar som
kulturplatser ställs inför och identifiera god praxis.
Vi hoppas att revisionen ska bidra till kunskap om relevansen och
ändamålsenligheten hos EU:s insatser för kulturplatser. På ett mer allmänt plan är vår
tanke att den också ska bidra till den pågående debatten om kulturens plats i EU.
Iakttagelser
Den befintliga ramen för EU:s investeringar i kulturplatser
saknar fokus, och samordningen är begränsad
Den strategiska ramen för EU:s insatser för kultur är komplex och
återspeglas endast delvis i EU:s finansiering
En lämplig ram för EU:s investeringar i kulturplatser är av central betydelse för att
maximera investeringarnas effekter när det gäller att uppnå de mål som fastställts i
ramen. En förutsättning för det är en tydlig strategisk ram för EU:s insatser på
kulturområdet, med en stark samordning mellan den rättsliga ramen (dvs.
lagstiftningen om EU:s fonder) och den icke-rättsliga ramen (dvs. strategier). Mål bör
fastställas tydligt utifrån identifierade behov och åtgärder utformas på motsvarande
sätt. Målen bör vara realistiska och uppnås genom lämpliga politiska instrument och
lämplig finansiering. Kraven på intressenter bör fastställas i överensstämmelse med
deras behörighet. För att framstegen mot måluppfyllelse ska kunna bedömas är det en
grundförutsättning att ramen övervakas.
Flera olika strategiska EU-ramar förekommer samtidigt, vilket påverkar EU:s insatser
på kulturområdet
EU:s strategiska inriktning har formulerats i tioårsplaner (Lissabonstrategin och
Europa 2020-strategin). Dessa planer behandlar inte kultur och är inte heller
synkroniserade med kommissionens femåriga mandatperiod eller med EU:s sjuåriga
finansieringsperioder.
Vad beträffar utformningen av kulturpolitiken på EU-nivå har EU infört en ram
som omfattar flera ansvarsnivåer (se punkterna 04–07). På den högsta nivån definieras
ramen av fördragen och EU:s internationella åtaganden (t.ex. Unescos konvention om
skydd för och främjande av mångfalden av kulturyttringar från 2005). Den preciseras i
kommissionens agendor och rådets fyraåriga arbetsplaner för kultur som tillsammans
bildar EU:s centrala ram för kultur. Flera dokument av strategisk betydelse
kompletterar ramen (se bilaga VI). I en tidigare publikation rapporterade vi att det
faktum att det finns flera strategiska ramar med överlappande perioder och mål är
komplext och kan vara förvirrande (se bild 1)16.
Punkterna 16–18 i revisionsrättens briefingdokument om en prestationsinriktad
sammanhållningspolitik, juni 2019.
Utgifter
Lissabonfördraget 2007
Maastrichtfördraget 1992
Unescos konvention från 2005
2030-agendan för hållbar utveckling
Lissabonstrategin
Prodi-kommissionen
Europa 2020
Första Barroso-kommissionen
Andra Barrosokommissionen
Juncker-kommissionen
Kommissionen: agendor för kultur
EU:s
kulturstrategi
Internationella
EU:s
prioriteringar åtaganden
EUfördrag
Bild 1 – Tidslinje för händelser
Europeisk agenda för en kultur i en alltmer globaliserad värld
Rådet: arbetsplaner för kultur
2008–2010
Fleråriga budgetramen 2000–2006
2002 2003 2004 2005 2006
2011–2014
Fleråriga budgetramen 2007–2013
En ny europeisk agenda
för kultur
2015–2018
2019–2022
Fleråriga budgetramen 2014–2020
2021–2027
2009 2010 2011 2012 2013 2014 2015 2016 2017 2018 2019 2020 2021 2022
Källa: Revisionsrätten.
Komplexiteten förvärras av den parallella förekomsten av olika aktörer
(kommissionen, rådet och medlemsstaterna) som samtidigt utarbetar och genomför
insatser på kulturområdet utan systematisk hänvisning till kommissionens agendor.
Inom kommissionen beaktas (”integreras”) kulturella aspekter på en rad olika
politikområden, med olika ansvariga avdelningar.
Övervakningen av målen i kommissionens agenda för kultur är inte tillräckligt
utvecklad
De viktigaste gemensamma strategiska mål som vägleder EU:s insatser på
kulturområdet fastställs i kommissionens agendor (se punkt 06). De omvandlas inte till
tydliga operativa mål. Trots att det finns många exempel på EU-åtgärder inom varje
mål, är det oklart vad EU försöker uppnå genom dessa åtgärder. Den nya agendan
innehåller varken bestämmelser om övervakning av hur de fastställda målen uppfylls
eller indikatorer för att mäta framsteg. Enligt kommissionen beror detta på att
kommissionen och medlemsstaterna inte har gemensamt fastställda mål, indikatorer
eller målvärden för utformningen av kulturpolitiken. Kommissionen använder sig inte
heller av de indikatorer som finns tillgängliga på programnivå, det vill säga de
indikatorer som fastställts i de olika EU-programmen, för att bedöma hur
framgångsrikt den nya agendan genomförs.
Inom ramen för rådets arbetsplaner för kultur vidtas samordnade åtgärder med
medlemsstaterna på detta område genom en icke bindande, mellanstatlig ram för
samarbete mellan medlemsstater som kallas den öppna samordningsmetoden. Enligt
kommissionen ”återstår utmaningen att föra över [den öppna samordningsmetodens]
rekommendationer till beslutsfattandet på nationell och europeisk nivå” 17. Även om
de kulturpolitiska ramar som medlemsstaterna i vårt urval hade infört i stort sett följde
de ekonomiska och sociala målen i den nya agendan, hänvisade ingen specifikt till den
nya agendan, och endast två hänvisade till 2007 års agenda.
Kommissionens agenda beaktas inte i de viktigaste EU-fonder som tillhandahåller
finansiering till kultur
När det gäller EU-finansiering är kultur i första hand ett medel att uppnå andra
EU-prioriteringar och mål (t.ex. stödja stadsutveckling och regional utveckling,
företagande och turism) och inte i sig en huvudprioritering. Dessa prioriteringar
hanteras genom andra EU-fonder. Den enda EU-fond som har utformats för kultur är
programmet Kreativa Europa, men det är väldigt litet sett till finansieringen. Det
fördelar runt 209 miljoner euro per år från EU-budgeten 18 till kultur i 28
medlemsstater och åtta länder utanför EU. Det beloppet motsvarar de årliga
driftskostnaderna för vissa enskilda kulturplatser. Till exempel uppgick Parisoperans
kostnader till 200,8 miljoner euro 2018 19.
Av de tolv EU-fonder som potentiellt skulle kunna stödja kultur som vi
analyserade hänvisar endast förordningen om Kreativa Europa till kommissionens
agenda från 2007 (se bilaga II). De två på varandra följande agendorna från
kommissionen fastställdes efter det att de fleråriga budgetramarna för ESI-fonderna
hade införts (se bild 1) och kunde därför inte beaktas i ESI-fonderna.
Kommissionen har utvecklat flera initiativ som kan främja kulturplatser,
men samordningen med finansieringsarrangemang är begränsad
En lämplig ram för EU:s investeringar i kulturplatser behöver ha ändamålsenliga
arrangemang för samordning mellan de olika politikområden som bidrar till främjandet
av kulturplatser. Samordnade åtgärder inom kommissionen kan säkerställa
Kommissionens rapport om genomförandet och betydelsen av arbetsplanen för kultur
2011–2014, COM(2014) 535 final, 25.8.2014, s. 12, och kommissionens rapport om
genomförandet av den europeiska kulturagendan, COM(2010) 390 final, 19.7.2010, s. 8.
Se artikel 24 i programmet Kreativa Europa.
Årlig prestationsöversyn – kulturutgifter, bilaga till lagförslaget om ansvarsfrihet, Frankrikes
finansministerium, 2018, s. 223.
komplementaritet mellan EU-fonder och garantera en effektiv användning av de
ekonomiska resurserna så att de föreslagna initiativen kan utvecklas.
Kommissionen har utvecklat flera initiativ som syftar till att främja kulturplatser
Kommissionen har det senaste årtiondet tagit fram en lång rad initiativ som syftar
till att främja kulturplatser, särskilt på kulturarvsområdet. Det senaste av dem är
Europaåret för kulturarv 2018, som resulterade i en europeisk ram för insatser för
kulturarvet 20 och som var den första europeiska sektorsövergripande och integrerade
kulturarvsstrategin. Exempel på andra initiativ är priser och utmärkelser för att främja
hållbar turism eller uppmärksamma en viss kulturplats (se tabell 2).
Tabell 2 – EU-märkningar och EU-priser för att främja kulturplatser
Utmärkelse/Pris
Beskrivning
Europeiska kulturhuvudstäder
(sedan 1985)
Två olika europeiska städer utses årligen till europeiska
kulturhuvudstäder i syfte att lyfta fram deras kulturliv
och kulturella utveckling.
EU:s kulturarvspris
(sedan 2002)
Främjar bästa praxis när det gäller bevarande av
kulturarvet, förvaltning, forskning, utbildning och
kommunikation.
Framstående europeiska
resmål (sedan 2006)
Främjar hållbar turism genom att öka synligheten för nya,
icke-traditionella europeiska destinationer.
Europeiska kulturarvsmärket
(sedan 2013)
Tilldelas kulturarvsplatser som har ett symboliskt
europeiskt värde. Det omfattar även det immateriella
kulturarvet.
Logotypen för Europaåret för
kulturarv (sedan 2018)
Logotyp som används under de evenemang och
festligheter som anordnas i samband med Europaåret för
kulturarv.
Europeisk huvudstad för smart
turism (sedan 2019)
Belönar turistmål för deras hållbarhet, tillgänglighet,
digitalisering, kulturarv och kreativitet.
Källa: Revisionsrätten.
Myndigheterna i de medlemsstater som vi besökte ansåg att initiativet
Europeiska kulturhuvudstäder var särskilt gynnsamt (i ruta 1 ges exempel på positiva
effekter som de portugisiska myndigheterna beskrev för oss). En av de granskade
stödmottagarna bekräftade att den hade noterat en betydande ökning av antalet
besökare när Wrocław var europeisk kulturhuvudstad 2016. De experter vi intervjuade
Arbetsdokument från kommissionens avdelningar, SWD(2018) 491, 5.12.2018.
lovordade även några av kommissionens nyare initiativ (t.ex. Europaåret för kulturarv
och den nya agendan).
Ruta 1
Exempel på positiva effekter av initiativet Europeiska
kulturhuvudstäder
Guimarães i Portugal var europeisk kulturhuvudstad 2012. Enligt den studie som
medlemsstatens myndigheter gjorde i efterhand omfattade initiativet
investeringar i kulturell infrastruktur och stadsförnyelse på omkring 41,7 miljoner
euro i stödberättigande kostnader samt ett kulturprogram som genomfördes
under hela 2012. Under samma år uppskattas antalet övernattningar i regionen ha
ökat med 43 %, vilket skapade 2 111 jobb.
Invigning av Guimarães som europeisk kulturhuvudstad
© Capital Europeia da Cultura Guimarães 2012.
Källa: Interimsrapport om de sociala och ekonomiska effekterna av Guimarães 2012.
På internationell nivå kan kulturplatser få andra utmärkelser (se bilaga VII). Den
samtidiga förekomsten av flera olika utmärkelser och priser gör att det är svårt att
tydligt avgöra vilket värde de är tänkta att tillföra.
Samordningen av kommissionens kulturinitiativ med Erufs finansieringsarrangemang
är begränsad
Vi analyserade hur GD Utbildning, ungdom, idrott och kulturs kulturinitiativ hade
samordnats med Eruf. Framför allt frågade vi stödmottagarna i de besökta projekten
vilka effekter Europeiska kulturarvsmärket och andra kommissionsinitiativ hade haft.
Kommissionens kulturinitiativ har mycket begränsad effekt på stödmottagares tillgång
till Eruf-medel. Varken Eruf-förordningen eller de operativa program inom Eruf som
omfattades av revisionen innehåller bestämmelser som gagnar projekt som redan
deltar i ett av kommissionens kulturinitiativ.
Finansieringsarrangemang finns tillgängliga för Unescos världsarvsplatser inom
Eruf. För programperioden 2014–2020 fastställer den nuvarande Eruf-förordningen ett
högre tak för Unescos världsarvsplatser (maximalt 20 miljoner euro i Erufmedfinansieringsstöd till Unescos världsarvsplatser och 10 miljoner euro till andra
kulturplatser)21. Unesco-utmärkelsen användes också som kriterium för att välja ut
projekt i fem av de 21 urvalsförfaranden som vi granskade. Myndigheterna i
medlemsstaterna ansåg även att nationella utmärkelser var viktiga, och i fyra av de
granskade urvalsförfarandena gynnades projekt med sådana utmärkelser.
Vårt urval av projekt innehöll två platser som fått Europeiska kulturarvsmärket
och en plats som deltog i initiativet Europeiska kulturhuvudstäder. När myndigheterna
i medlemsstaterna valde ut projekt för Eruf-finansiering betraktades inte kulturplatsers
deltagande i EU-initiativ som ett kriterium (se bilaga V). Detta föreslog inte heller
kommissionen i sina kommentarer innan den godkände de operativa programmen.
Den europeiska panel som ansvarar för övervakningen av europeiska kulturarvsplatser
har angett att brist på finansiering till platser som fått utmärkelsen skulle kunna
äventyra utmärkelsens hållbarhet och synlighet 22. Utmärkelsen är också en
angelägenhet för parlamentet, som har rekommenderat att den ges större synlighet 23.
Komplementariteten mellan EU-fonder är inte tillräckligt synlig när det gäller
investeringar i kulturplatser
I enlighet med principen om integrering är genomförandet av de mål som
fastställts i kommissionens agenda från 2007 i praktiken utspritt på olika
politikområden och får stöd genom olika fonder som förvaltas av 15 olika
generaldirektorat inom kommissionen. Samordningen mellan de olika direktoraten
sker huvudsakligen genom en avdelningsövergripande arbetsgrupp för kultur och
kulturarv och genom samråd mellan avdelningar när program och förordningar ska
antas.
Artikel 3.1 i förordning (EU) nr 1301/2013 om Eruf, ändrad genom förordning (EU, Euratom)
2018/1046 av den 18 juli 2018 om finansiella regler för unionens allmänna budget (EUT
L 193, 30.7.2018, s. 1).
Panel Report on Monitoring, Europeiska kulturarvsmärket, 19 december 2016.
Europaparlamentets resolution av den 2 mars 2017 om genomförande av programmet
Kreativa Europa, P8_TA(2017)0062.
Resultaten av den samordningen framgår inte tydligt i de olika EU-
fondförordningarna. Även om förordningarna i olika grad speglar vissa delar av
agendan från 2007, hänvisar inte någon av dem (utom den som gäller Kreativa Europa)
specifikt till den, och merparten av dem har inte kultur som mål (se punkt 24 och
bilaga II).
I förordningen om gemensamma bestämmelser24 föreskrivs arrangemang för att
främja samordning mellan fonder genom att det införs en gemensam strategisk ram
och ett krav att medlemsstaterna ska rapportera om arrangemangen för samordning
mellan EU-fonder i partnerskapsöverenskommelserna och de operativa programmen.
Särskilt när det gällde kulturplatser identifierade vi brister i dessa
samordningsarrangemang.
För det första: Även om kulturarvsplatser potentiellt kan finansieras genom olika
ESI-fonder beroende på vilka mål de har, bedömer kommissionen inte
komplementaritet och möjliga synergieffekter i användningen av EU-fonder specifikt
för kulturarvsplatser när den antar partneröverenskommelser och operativa program.
De samordningsarrangemang som beskrivs i partnerskapsöverenskommelserna och de
operativa programmen är allmänna och hänvisar inte alltid specifikt till kulturplatser.
Vi analyserade särskilt hur Ejflu-investeringar i kulturplatser hade särskilts från Erufinvesteringar i kulturplatser i partnerskapsöverenskommelserna, de nationella Ejfluprogrammen och de operativa programmen inom Eruf. I fyra medlemsstater var
skillnaderna oklara mellan de två fonderna, som potentiellt skulle kunna finansiera
samma typ av projekt.
För det andra nämndes inte samordning med Kreativa Europa eller dess
föregångarfond (”programmet Kultur” 25) i urvalet av strategiska dokument från tre
medlemsstater som ingick i revisionen. På projektnivå, för det tredje och slutligen,
belönade fyra av de 21 bedömda urvalsförfarandena i vårt urval specifikt
komplementaritet med andra EU-fonder som ett kriterium för finansiering, dock utan
att Kreativa Europa nämndes särskilt. Detta fick till följd att ett projekt inom Kreativa
Europa kompletterade ett Eruf-projekt på endast en av kulturplatserna i vårt urval.
Förordning (EU) nr 1303/2013 om allmänna bestämmelser för ESI-fonderna (EUT L 347,
2013, s. 320).
Beslut nr 1855/2006/EG av den 12 december 2006 om inrättande av programmet Kultur
(2007–2013) (EUT L 372, 27.12.2006, s. 1).
Eruf är ett instrument för att strukturera medlemsstaternas
investeringar i kulturplatser, men sådana investeringar behandlas inte
som en prioritering för Eruf
I en lämplig ram för investeringar i kulturplatser bör de EU-fonder med mest
finansiering tillgänglig för sådana investeringar, särskilt Eruf, spegla EU:s kulturella ram
i sina åtgärder. För det ändamålet bör kommissionens mål på kulturområdet tydligt
återspeglas i medlemsstaternas partnerskapsöverenskommelser och operativa
program.
EU:s totala utgifter för investeringar i kulturplatser övervakas inte specifikt
Även om utgifterna för kultur endast utgör en liten del av den samlade Eruf-
budgeten (runt 4,7 miljarder euro har planerats för programperioden 2014–2020, eller
2,3 %), är Eruf den viktigaste källan till EU-finansiering av investeringar i kulturplatser.
Enligt förordningen om gemensamma bestämmelser ska myndigheterna i
medlemsstaterna rapportera utgifter per insatskategori. En sådan är ”Skydd, utveckling
och främjande av offentliga kulturtillgångar och kulturarv”. Men kategorin är bredare
än infrastrukturinvesteringar, och medlemsstaterna använder den inte på samma sätt.
I bilaga VIII presenteras hur omfattningen av Erufs investeringar i kultur har utvecklats
och övervakningsarrangemangen för dem.
År 2014 gjorde kommissionen en kartläggning av tillgängliga EU-medel för
kulturarvsinsatser 26. Kartläggningen var inte uttömmande 27. Den innehöll inga
detaljerade och aktuella uppgifter om vilka EU-belopp som anslagits och använts till
kulturarvsinsatser, inbegripet tillhörande fysiska investeringar. Dessa uppgifter är inte
kända eftersom inte alla olika EU-fonder kräver att medlemsstaterna och
stödmottagarna systematiskt lämnar information om kulturåtgärder.
Kommissionen har försökt harmonisera olika typer av statistiska data om
offentliga utgifter för kultur och deras effekter. Den grundläggande referensen för EU:s
kulturstatistik är en rapport från det europeiska statistiska systemnätet för kultur från
Mapping of Cultural Heritage actions in the European Union policies, programmes and
activities, 2014 års version (https://www.europa-creativa.eu/Files/uploads/29-2014heritage-mapping_en.pdf) och en uppdaterad version från 2017
(https://ec.europa.eu/culture/sites/culture/files/2014-heritage-mapping-version2017_en.pdf).
Mapping of Cultural Heritage actions in the European Union policies, programmes and
activities, versionerna från 2014 och 2017, s. 2.
Eurostat har följt upp nätets arbete 29. Att stärka evidensbasen på EU-nivå är
också en av huvudprinciperna för den nuvarande europeiska ramen för åtgärder för
kulturarv20. Men än så länge finns det ingen obligatorisk EU-ram för insamling av data
och rapportering om kultur eller kulturplatser.
Eruf tillhandahåller en ram för medlemsstaternas investeringar i kulturplatser
I en granskningsrapport från 201730 konstaterade vi att den nuvarande Eruf-
förordningen föreskriver ett mer strukturerat tillvägagångssätt för EU-insatser jämfört
med programperioden 2007–2013 genom att den kräver att de operativa programmen
tydligare ska ange insatsernas mål (särskilda mål/resultat) och hur de förväntas uppnås
(nödvändig finansiering, åtgärder som ska vidtas och förväntad output). Detta gäller
särskilt när åtgärder utformas efter investeringsprioriteringar, såsom kulturarv
(se punkt 44).
Ramen för 2014–2020 har också förbättrats när det gäller indikatorer för att mäta
Erufs stöd till kulturplatser, och den nuvarande förordningen fastställer en gemensam
outputindikator avseende kulturplatser. Till programperioden 2021–2027 föreslår
kommissionen att antalet gemensamma indikatorer avseende kulturplatser ska ökas
och, för första gången, att gemensamma resultatindikatorer ska tas med
(se bilaga VIII). I ett yttrande nyligen välkomnade vi införandet av gemensamma
indikatorer och konstaterade att de är ett viktigt steg mot en ökad inriktning på
resultat och prestation 31.
Eruf-ramens betydelse framgår av de tre besökta medlemsstaternas
kulturstrategier. I Polens kulturstrategi betraktas kultur som ett medel att uppnå den
ekonomiska och sociala sammanhållning som eftersträvas av Eruf. I Italien har
regeringen tagit fram ett nationellt finansieringsprogram som ska komplettera det
nationella operativa programmet för kultur inom Eruf 32 med samma mål och
finansieringskriterier. I Portugal begärde kommissionen att en kartläggning skulle göras
av EU-finansieringen där behoven av investeringar i kulturplatser analyserades och
investeringsprioriteringar identifierades.
Final Report of the European Statistical System Network on Culture (ESSnet-Culture), 2012.
Se t.ex. Guide to culture statistics, Eurostat, 2018 års upplaga.
Särskild rapport 02/2017 Kommissionens förhandlingar om partnerskapsöverenskommelser
och program inom sammanhållningspolitiken 2014–2020: utgifterna riktas mer mot Europa
2020-prioriteringar, men arrangemangen för resultatmätning är allt mer komplexa.
Punkt 59 i revisionsrättens yttrande nr 6/2018.
Programma di Azione e Coesione Complementare al PON Cultura e Sviluppo 2014–2020.
Eruf är en viktig källa till finansiering av offentliga investeringar i kulturplatser i vissa
medlemsstater
Eruf-förordningen fastställer en rad tematiska mål och investeringsprioriteringar
som medlemsstaterna kan välja beroende på vilka behov de har. Under
programperioden 2014–2020 avser stödet till kulturplatser specifikt kulturarvsplatser
inom investeringsprioritering 6 c ”bevara, skydda, främja och utveckla natur- och
kulturarvet” inom det tematiska målet ”att bevara och skydda miljön och främja en
hållbar användning av resurser”. Kulturplatser kan också stödjas inom andra
investeringsprioriteringar, nämligen genom Erufs stöd till innovation (tematiskt mål 1)
eller små och medelstora företags konkurrenskraft (tematiskt mål 3) eller när de ingår i
en bredare territoriell utvecklingsstrategi som främjar sysselsättning (tematiskt mål 8)
eller social delaktighet (tematiskt mål 9). Stadsförnyelse, inom investeringsprioritering
e, är också en vanlig prioritering som väljs ut i de operativa programmen för att
stödja kulturplatser.
Under perioden 2010–2017 uppgick investeringarna i kulturplatser med Eruf-
medel till cirka 750 miljoner euro per år. De stod för över 25 % av alla offentliga
investeringar i kulturella tjänster i runt en tredjedel av medlemsstaterna och för över
% i Portugal och Grekland (se figur 1). Fonden var därför en viktig källa till
finansiering av investeringar i kulturplatser i många medlemsstater. På projektnivå
skulle, enligt vår enkät, 44 % av projekten inte ha genomförts utan Eruf-stöd, och 48 %
skulle ha skjutits upp eller genomförts i reducerad omfattning.
Figur 1 – Eruf-finansiering och medlemsstaternas kapitalinvesteringar i
kulturplatser, årligt genomsnitt 2010–2017
miljoner euro
1 000
1 500
2 000
2 500
3 000
3 500
Grekland
Portugal
57,8 %
Cypern
49,8 %
Malta
46,9 %
Bulgarien
37,8 %
Litauen
35,3 %
Rumänien
28,7 %
Slovenien
28,3 %
Slovakien
26,1 %
Ungern
22,2 %
Polen
21,9 %
Tjeckien
21,3 %
Kroatien*
18,2 %
Lettland
9,2 %
Italien
9,2 %
Estland
7,1 %
Genomsnitt EU-28
6,8 %
Spanien
Offentliga investeringar i
kulturella tjänster (årligt
genomsnitt 2010–2017)
% av Erufs finansiering som gått
till kulturplatser (årligt
genomsnitt 2010–2018)
5,4 %
Tyskland
2,3 %
Belgien
2,2 %
Finland
1,6 %
Nederländerna
1,3 %
Förenade kungariket
1,0 %
Danmark
0,7 %
Frankrike
0,6 %
Sverige
0,6 %
Österrike
0,4 %
Luxemburg
0,0 %
Irland
0,0 %
Anm.: 1) Vi har använt Eurostats data om offentliga utgifter för kulturella tjänster (COFOG: GF08.2) för
att uppskatta medlemsstaternas investeringar i kulturplatser. Detta är den bästa uppskattning som finns
tillgänglig. Kapitalinvesteringar i kulturella tjänster inbegriper: investeringsbidrag (D92), fasta
bruttoinvesteringar (P.51g) och anskaffning minus avyttringar av icke finansiella icke producerade
tillgångar (NP). Siffrorna representerar ett årligt genomsnitt av de belopp som använts av nationella och
lokala myndigheter (offentliga utgifter) under åren 2010–2017. 2) Eruf-investeringar i kulturplatser,
uttryckt som ett årligt genomsnitt, inkluderar de utgifter som bokförts för kulturplatser under
programperioderna 2007–2013 och 2014–2020 (fram till 2018).
* När det gäller Kroatien har endast medel som använts under den nuvarande programperioden
beaktats.
Källa: Revisionsrätten, på grundval av Eurostat, General government expenditure by function (COFOG),
onlinedatakod: [gov_10a_exp], plattformen för öppna data om sammanhållningspolitiken och
kommissionens information.
På nationell nivå fann vi exempel på hur medlemsstater diversifierar
inkomstkällorna för kulturplatser och utvecklar finansieringssystem som bygger på
privata medel (se ruta 2). Diversifiering av finansieringen av kulturarvet är även ett av
de ämnen som rådet behandlar i arbetsplanen för kultur 2019–2022 33.
Ruta 2
Exempel på finansieringssystem som tagits fram på nationell nivå
Kulturarvslotteri (Frankrike): Med Förenade kungariket som förebild införde den
franska regeringen ett nationellt kulturarvslotteri 2018 för att stödja
restaureringen av några ikoniska lokala kulturarvsplatser (20 miljoner euro
samlades in det året till restaureringen av 18 platser).
Kulturarvslotteri (Italien): Sedan 1997 reserveras en del av lotteriintäkterna för
ministeriet med ansvar för kulturarvet och fördelas till en lång rad
kulturarvsprojekt i hela Italien som avser återställande och bevarande av
kulturarvet, inbegripet arkeologiska, historiska, konstnärliga och arkiv- och
biblioteksrelaterade projekt samt till återställande av landskapsarkitektur och
kulturella verksamheter. Ett projekt i vårt urval, Ex-Convento di Sant’ Antonio, fick
omkring 2,4 miljoner euro från ”Programma Triennale Lotto 2007–2009”. Panteon
i Rom och den grekiska teatern i Syrakusa är andra exempel på kulturplatser som
finansierats.
Korrigerande beskattning (Polen): Polen inrättade en ny fond 2018 för att
finansiera skydd och renovering av historiska platser. Finansieringen kommer från
de administrativa böter som utdöms för överträdelser av kraven på skydd av
historiska platser.
Investeringar i kulturplatser behandlas inte som en prioritering för Eruf
Eruf syftar till att främja ekonomisk, social och territoriell sammanhållning, som
är en av EU:s viktigaste uppgifter enligt EU-fördraget 34. Denna uppgift har tillsammans
med målen för Europa 2020-strategin om smart och hållbar tillväxt för alla lett till att
Erufs ram är centrerad kring ekonomiska och sociala överväganden. Investeringar i
kulturplatser är därför ett medel att uppnå ett mål och ska finansieras endast om de
har en socioekonomisk effekt.
Se punkt Error! Reference source not found..
Artikel 3.3 i EU-fördraget.
Utöver denna socioekonomiska grund infördes genom Eruf-förordningen 2014–
restriktioner för Erufs investeringar i kulturplatser som innebär att endast
småskalig infrastruktur finansieras. Det är oklart hur denna bestämmelse bidrar till de
mål som fastställts i kommissionens agendor för kultur. I den ursprungliga
förordningen framgick det inte heller klart vad som avsågs med ”småskalig”, vilket
skapade osäkerhet kring vilka typer av projekt Eruf kunde finansiera.
Olika tolkningar gjordes av Eruf-restriktionen. Först definierade kommissionen
småskalig” administrativt som investeringar på upp till 5 miljoner euro (10 miljoner
euro för Unescos världsarvsplatser)35. Efter det att elva medlemsstater hade framfört
ett klagomål till kommissionen 36 uppgav kommissionen att flexibilitet kunde tillämpas
när det gällde hur olika småskaliga infrastrukturobjekt kunde få stöd inom en enda
integrerad insats. Först fyra år senare förtydligade den ändrade Eruf-förordningen för
2014–2020 den rättsliga grunden och fastställde taket för berättigande av Eruf-stöd till
miljoner euro (20 miljoner euro för Unescos världsarvsplatser).
På grund av denna finansieringsrestriktion granskade kommissionen investeringar
i kulturplatser under förhandlingarna om 2014–2020, och investeringarna var inte en
prioritering inom Eruf. I de tre besökta medlemsstaterna, och när det gällde de
operativa programmen och partnerskapsöverenskommelserna i vårt urval, hade
kommissionen inte identifierat investeringar i kultur som ett prioriterat område under
förhandlingarna utan framfört ståndpunkten att kultur endast skulle behandlas genom
e-kultur 37 (Italien och Polen) och i samband med främjande av kulturella och kreativa
näringar 38 (Polen och Portugal). Kommissionen föreslog även en minskning av anslagen
till kulturella investeringar (Polen och Italien) och införde finansieringsrestriktioner i
samtliga fall.
Medlemsstaternas kulturpolitik bedöms inte specifikt inom Eruf. När det gäller
partnerskapsöverenskommelserna och de operativa programmen i vårt urval krävde
inte kommissionen att medlemsstaterna skulle planera kulturinsatserna i
överensstämmelse med kommissionens europeiska agenda för kultur när den antog
dem för programperioden 2014–2020.
Kommissionens avdelningar, riktlinjer för handläggare, definition av ”småskalig” när det
gäller infrastruktur enligt Eruf-förordningen, version 1.0, 7 juli 2014.
Informerande not från den polska delegationen till rådet, The necessity of raising the
maximum value of small-scale cultural infrastructure implemented within the European
Regional Development Fund 2014–2020, 8561/15, 6 maj 2015.
Inom tematiskt mål 2 ”Att öka tillgången till, användningen av och kvaliteten på IKT”.
Inom tematiskt mål 3 ”Att öka konkurrenskraften för SMF”.
Varierande ändamålsenlighet och hållbarhet hos de granskade
Eruf-projekten
Vi bedömde ändamålsenligheten i Eruf-projekt avseende kulturplatser baserat på
hur projektens mål och planerade resultat hade uppnåtts. Framför allt bedömde vi hur
de ekonomiska, sociala och kulturella målen hade uppfyllts. Genomförandet av dessa
mål skapar externa effekter i samhället.
Vi bedömde hållbarhet som platsens förmåga att fortsätta verksamheten, vilket
kräver regelbundet underhåll och, vid behov, restaurering av den fysiska
infrastrukturen. Det krävs också tillgång till ekonomiska och personella resurser. Detta
handlar om kulturplatsernas interna verksamhet.
De beskrivna målen och hållbarhetsfaktorerna är sammanlänkade (se bild 2). I
princip har ett kulturinvesteringsprojekt effekter på uppfyllelsen av alla tre målen och
på kulturplatsens hållbarhet. Effekterna kan emellertid ha motstridiga inriktningar.
Ekonomiska mål kan öka den ekonomiska hållbarheten för en plats men hindra
bevarandet av den (t.ex. överturism och minskade underhållskostnader). Vissa sociala
mål kan leda till minskande ekonomisk hållbarhet (t.ex. minskade inträdesavgifter)
eller hindra bevarandet av en plats (t.ex. för många besökare). Kulturella mål kan öka
den sociala delaktigheten och skapa ekonomiska effekter men kan också ha negativ
inverkan på platsens ekonomiska hållbarhet (t.ex. kostnadsökningar när utbudet av
kulturaktiviteter ökar).
Bild 2 – Samband mellan ändamålsenlighet och hållbarhet för
kulturplatser
Socialt mål
Hållbarhet
Kulturellt
mål
Restaurering
Och
underhåll
Resurser
Ekonomiskt
mål
Källa: Revisionsrätten.
De slutförda, granskade projekten var operativa, deras mål var för det
mesta ekonomiska och det gick inte alltid att säga om de hade uppnåtts
Eruf-projekten ska uppnå de mål som har fastställts vid projekturvalet. För att
mäta måluppfyllelsen ska stödmottagarna i Eruf-projekt fastställa relevanta indikatorer
och på ett tillförlitligt sätt rapportera hur målvärdena uppnås. När Eruf-projekten har
slutförts ska kulturplatserna vara i drift och bidra till uppfyllelsen av mål i de operativa
program som de får finansiering från.
De granskade operativa programmen och projekten inom Eruf var främst inriktade
på ekonomiska mål och mindre på sociala och kulturella mål
I enlighet med Eruf-målen använde alla operativa program i vårt urval
kulturplatser som en resurs för förbättring av ekonomins konkurrenskraft eller för
territoriell utveckling (se bilaga IX). Detta skedde genom främjande av turism eller
strategier för stadsutveckling (se ruta 3).
Ruta 3
Exempel på en strategi för stadsutveckling
Katowice är huvudstad i regionen Śląskie (Schlesien) och centrum i det största
stadsområdet i södra Polen med 4,8 miljoner invånare. Regionen blomstrade på
1800-talet tack vare den snabba utvecklingen av gruv- och stålindustrin. I slutet av
1990-talet inledde Katowice en strategisk omorientering och gjorde kultur till en
central prioritering för staden.
Det granskade projektet, Polens nationella radiosymfoniorkester (NOSPR), är ett
resultat av den strategin. Fram till 2006 var det område där NOSPR nu har sina
lokaler, i hjärtat av staden, en före detta kolgruva.
Före detta kolgruva i centrala Katowice i Polen
© Katowices stad.
Källa: Katowices stad.
Förutom NOSPR byggde staden under en tioårsperiod i samma område även ett
internationellt kongresscentrum och ett museum (Muzeum Śląskie w Katowicach).
De tre stora investeringarna uppgick till totalt cirka 231 miljoner euro och
genomfördes med omfattande Eruf-stöd (123 miljoner euro). För investeringarna
utsåg Unesco Katowice till ”kreativ musikstad” 2015, och 2018 stod Katowice värd
för FN:s klimattoppmöte.
Område efter upprustning i Katowice i Polen
© Katowices stad.
Källa: Katowices stad.
Ekonomiska måls företräde framgår när resultatindikatorerna inom operativa
program och på projektnivå bedöms. Vad beträffar de granskade insatsområdena
syftar 26 av de 32 fastställda resultatindikatorerna till att fånga upp Eruf-insatsernas
ekonomiska effekter. Bilaga IX sammanfattar hur de olika målen för de granskade
insatsområdena mäts genom resultatindikatorer. Den visar den ekonomiska
dimensionens betydelse och att alla granskade insatsområden har ett ekonomiskt mål
under båda programperioderna.
På projektnivå mäter alla resultatindikatorer som stödmottagarna valt ut i de
granskade projekten för perioden 2014–2020 och 45 av de 59 resultatindikatorerna för
programperioden 2007–2013 projektens ekonomiska effekter (se figur 2).
Figur 2 – Andel (antal) indikatorer i de granskade projekten som mäter
de kulturella, sociala och ekonomiska målen
% (12)
% (10)
% (45)
Ekonomiska
Sociala
% (25)
% avser antalet
besökare
% (11)
Kulturella
% avser
antalet besökare
% (0)
Resultatindikatorer för 2007–2013 Resultatindikatorer för 2014–2020
Anm.: 1) Under perioden 2014–2020 finns det endast fem projekt med resultatindikatorer. 2) Varje
indikator kan mäta mer än ett mål, varför summan kan vara högre än 100 %.
Källa: Revisionsrätten.
När det gäller sociala mål har kommissionens agendor, parlamentet39 och rådet40
ofta gett uttryck för att det är nödvändigt att stärka kulturinsatsernas sociala effekter.
Särskild uppmärksamhet har ägnats åt integrering av migranter, främjande av
jämställdhet mellan könen och arbete i partnerskap mellan kultursektorn och andra
sektorer. Vid ett informellt möte nyligen mellan EU-medlemsstaternas ministrar med
ansvar för Europafrågor och kulturministrar, om skydd av kulturarvet, pekades på
behovet av att främja den europeiska ungdomens engagemang för och medvetenhet
om kulturarvet 41.
Europaparlamentets resolution av den 2 mars 2017 om genomförande av programmet
Kreativa Europa, P8_TA(2017)0062, och förslag till Europaparlamentets
lagstiftningsresolution om förslaget till inrättande av programmet Kreativa Europa (2021–
2027), A8-0156/2019, 4.3.2019.
Rådets slutsatser om de kulturella och kreativa sektorernas samverkan med andra sektorer
för att stimulera innovation, ekonomisk hållbarhet och social delaktighet (EUT C 172,
2015, s. 13).
Gemensam förklaring som antogs vid det informella mötet mellan EU-medlemsstaternas
kulturministrar och ministrar med ansvar för Europafrågor om skydd av det europeiska
kulturarvet, Paris, 3 maj 2019.
De granskade insatsområdena med sociala mål syftar framför allt till att förbättra
kulturplatsers tillgänglighet eller öka den sociala sammanhållningen. Den indikator
som används oftast för att mäta projekts sociala aspekter är antal besökare
(se figur 2). Den effekt som kulturplatser har på besökare, såsom välbefinnande, stöd
till missgynnade grupper eller främjande av utbildningsinsatser, registreras sällan med
särskilda indikatorer. Social verksamhet genomfördes likväl, i olika grad, i 10 av de 11
slutförda projekt som vi besökte (se ruta 4).
Ruta 4
Exempel på sociala verksamheter som utvecklats på en kulturplats
San Carlo-teatern i Neapel i Italien är det äldsta operahuset i världen som ännu är i
bruk. Teatern är inte bara ett operahus utan även en plats där besökarna kan gå
på dansföreställningar och konserter, besöka utställningar och muséet eller gå på
guidad tur. Teatern har särskilt fokus på att locka ungdomar. Förutom en
balettskola driver kulturplatsen i partnerskap med en förening även ett
utbildningsprojekt som finansieras av Kreativa Europa. Projektet, som syftar till att
lära barn från tidig ålder att sjunga och tycka om opera, ska först utbilda lärare
genom en rad musikkurser och därefter ge dem stöd när de undervisar elever i
skolorna. När musikutbildningen är klar anordnas en föreställning på teatern för
lärare, elever och familjemedlemmar. Eleverna uppträder och sjunger på scen,
ackompanjerade av professionella sångare och av teaterns orkester, klädda i
kostymer som de har tillverkat själva.
Teatro di San Carlo i Neapel i Italien
© Fotograf: Luciano Romano.
Arkitekt: Giovanni Antonio Medrano.
Källa: Teatro di San Carlo.
Vad beträffar kulturella mål syftade de insatsområden som vi granskade framför
allt till att bevara kulturarv. Alla de granskade insatsområdena hade inte ett tydligt
fastställt kulturellt mål, och de som hade det hade i de flesta fall inte fastställt
resultatindikatorer för att mäta måluppfyllelsen (se bilaga IX). I nästan hälften av de
granskade förfarandena ansåg inte de förvaltande myndigheterna inom Eruf att
kulturella aspekter var relevanta när de valde ut projekt (se bilaga V).
Alla slutförda, granskade projekt var operativa vid tidpunkten för revisionen, men
projektens prestation kan ofta inte bedömas
Alla de elva slutförda projekt som vi besökte var operativa vid tidpunkten för
revisionen, och förvaltningsteamen på platserna var engagerade i och verkade för att
bevara och främja dem. För att bedöma hur ändamålsenligt projekten uppfyllde sina
målvärden analyserade vi uppfyllelsen av 71 resultatindikatorer som hade rapporterats
av stödmottagarna i de 17 slutförda projekt som hade resultatindikatorer i vårt urval
(se bilaga IV).
Mindre än en tredjedel av de granskade projekten hade uppnått alla de
fastställda målvärdena inom den angivna perioden. Om de övriga projektens
prestation går det inte att dra någon slutsats (se figur 3). Vid tidpunkten för revisionen
hade dock ytterligare tre projekt nått sina målvärden. Vi noterade emellertid flera
brister i valet och rapporteringen av indikatorer.
Figur 3 – Projektens prestation: antal slutförda projekt som uppnått
fastställda målvärden för resultatindikatorer
När projektet har slutförts
Projekt som det inte
går att dra en
slutsats om
(en del målvärden
uppnådda, vissa inte
uppnådda och andra
kan inte bedömas på
grund av att
information saknas)
Källa: Revisionsrätten.
Projekt som inte
uppnådde något
målvärde
Projekt som uppnådde
alla målvärden
Projekt utan
resultatindikatorer
Vad gäller valet av indikatorer konstaterar vi att sex projekt inte hade några
resultatindikatorer alls. Det innebär att uppfyllelsen av projektmål inte kan mätas
genom resultatindikatorer för omkring en fjärdedel av de slutförda projekten.
Dessutom kan 16 av de 71 resultatindikatorerna inte användas till att dra slutsatser om
projektens ändamålsenlighet eftersom de inte är relevanta för projektmålen.
Ytterligare tolv är i själva verket inte resultat- utan outputindikatorer.
Alla de elva besökta projekt som hade slutförts vid tidpunkten för revisionen
hade resultatindikatorer. Vi analyserade tillförlitligheten hos de resultat som
stödmottagarna hade rapporterat för dessa indikatorer och konstaterade att 18 av de
rapporterade resultaten inte var tillförlitliga på grund av att resultat hade beräknats
felaktigt, att det saknades bevis som bekräftade resultaten eller att beräkningar inte
kunde verifieras (se tabell 3).
Tabell 3 – Tillförlitlighet hos rapporterade resultat för indikatorerna
inom de besökta, slutförda projekten (antal indikatorer)
Resultatindikatorer
Varav antal besökare
Totalt
Tillförlitliga
Ej tillförlitliga
felaktig beräkning
brist på bevis
icke verifierbara
beräkningar
Varav
Källa: Revisionsrätten.
Antal besökare” var den indikator som användes mest av stödmottagarna i de
besökta projekten, men den är ofta otillförlitlig (se tabell 3). Endast i två av de nio
slutförda, besökta projekten med indikatorer för antal besökare kunde vi få det antal
som hade rapporterats till de förvaltande myndigheterna att stämma. Dessutom är
kopplingen mellan ökningen av antalet turister och den typ av arbeten som utförts inte
alltid synlig. På tre av de elva kulturarvsplatser som vi besökte hade insatserna
begränsats till delrestaureringar (t.ex. renovering av tak eller av särskilda rum), vilket
inte direkt eller uteslutande leder till en ökning av antalet turistbesök.
Uppfyllelsen av de operativa programmens mål är inte direkt beroende av enskilda
projekts prestation
Redan i en av våra tidigare rapporter konstaterade vi att Erufs resultatindikatorer
för 2014–2020 inte är specifikt relaterade till de insatser som finansieras av
programmet 42. De resultatindikatorer som har fastställts i de granskade operativa
programmen för båda programperioderna har dessutom för det mesta begränsad
förmåga att mäta framsteg mot uppfyllelse. Nästan hälften av de operativa
programmens resultatindikatorer påverkas inte direkt av Eruf-projektens specifika
resultat utan av externa faktorer (se ruta 5). När det gäller mer än hälften av de
resultatindikatorer som definierats på projektnivå har uppfyllelsen av de fastställda
målvärdena ingen direkt påverkan på de resultat som uppnås på operativ programnivå
eftersom de operativa programmen inte omfattar dessa indikatorer.
Ruta 5
Exempel på en resultatindikator som fastställts för det operativa
programmet som inte mäter de direkta effekterna av projekten
Det portugisiska operativa programmet 2014–2020 för den centrala regionen
syftar till att främja regionen som ett framstående resmål. Detta sker genom
bevarande och turismfrämjande av kultur- och naturarvet. Eruf finansierar därför
renoverings- och restaureringsarbeten på kulturplatser, inklusive Unescos
världsarvsplatser.
För att mäta hur framgångsrika åtgärderna är innehåller det operativa
programmet resultatindikatorn ”antal övernattningar på hotell och andra
turistanläggningar i regionen”. År 2017 hade målvärdet för 2023 redan
överträffats med omkring 24 %, åtminstone delvis tack vare en turistboom i
medlemsstaten. Även om Eruf-projekten kan ha bidragit till detta resultat bör det
noteras att projekten bara hade börjat genomföras 2017 (inom insatsområde 7
hade åtaganden ingåtts för endast 68 % av de tillgängliga, totala, stödberättigande
kostnaderna). Eruf-projektens bidrag är därför begränsat och påverkas av externa
faktorer. Resultatindikatorn mäter inverkan av Erufs insatser snarare än
resultaten, det vill säga de direkta effekterna.
Punkterna 116 och 117 i revisionsrättens särskilda rapport 02/2017 Kommissionens
förhandlingar om partnerskapsöverenskommelser och program inom
sammanhållningspolitiken 2014–2020: utgifterna riktas mer mot Europa 2020prioriteringar, men arrangemangen för resultatmätning är allt mer komplexa.
Otillräcklig uppmärksamhet ägnas åt kulturplatsers hållbarhet
EU-investeringarnas hållbarhet måste säkerställas i alla faser av projektet. Det
första steget är att kontrollera, på ansökningsstadiet, att stödmottagarna har kapacitet
att driva eller fortsätta driva platsen. Därför bör kulturplatser som gagnas av EUinvesteringar ha ambitionen att bli självfinansierande i så stor utsträckning som
möjligt 43 (dvs. att deras verksamhetsintäkter täcker deras driftskostnader). Underhåll
är av grundläggande betydelse för bevarandet av kulturplatser och bör planeras
ordentligt för att begränsa kostnaderna för framtida arbeten och se till att platsens
skick inte försämras. Övervakningsarrangemang ska finnas på plats för att man ska
kunna bedöma om EU-investeringarna ger bestående resultat.
Inga Eruf-krav gäller bevarandet av kulturplatser som fått finansiering
Särskilt kulturarvsplatser behöver konstant underhåll och löper flera olika
bevaranderisker
Betydelsen av regelbundet underhåll för att kulturarvet ska bevaras slås fast i
Venedigdokumentet och Krakowstadgan 44. Alla stödmottagare som vi besökte
rapporterade att de regelbundet bedömer den fysiska statusen på sina kulturplatser,
men beslut om underhållsarrangemang fattas av stödmottagarna och kan ta sig olika
uttryck. ICOMOS har framhållit att kulturplatser i EU inte fokuserar tillräckligt på
förebyggande och regelbundet underhåll. Bara en besökt kulturplats hade en
uppdaterad, prioriterad och budgeterad flerårig underhållsplan. Det är god praxis och
ett krav för platser på Unescos världsarvslista 45 (se ruta 6) och rekommenderas för alla
kulturarvsplatser 46.
Kommissionens förslag till tematiska riktlinjer för handläggare om stöd till kultur-, turismoch idrottsrelaterade investeringar, version 1 – 13.5.2013.
Venedigdokumentet, internationell stadga för bevarande och restaurering av monument
och platser, 1964, och Krakowstadgan om principer för bevarande och restaurering av
byggnadsarvet, 2000.
Management Guidelines for World Heritage Sites, ICCROM, Unesco, ICOMOS, 1998 och
ICOMOS, Evaluations of Nominations of Cultural and Mixed Properties, Report for the World
Heritage Committee, 43rd session, WHC-19/43.COM/INF.8B1, 2019.
Artikel 4 i Venedigdokumentet.
Ruta 6
Exempel på en underhållsplan
Sedan 2015 har den arkeologiska parken i Pompeji en omfattande övervakningsoch underhållsplan för att skydda sina byggnader, sin konst och sina artefakter
från att förstöras. Planen består av olika delar och fastställer i) prioriterade
insatser som behövs för att bevara platsen med tillhörande tidsplan, ii) åtgärder
för att förbättra villkoren för parkens användning och för att främja turism, iii)
åtgärder för att minska riskerna för naturkatastrofer, iv) styrningsarrangemang
och v) övervakningsarrangemang. Sedan 2015 har platsen även ett digitalt arkiv
med information om utfört underhåll och efterföljande inspektioner.
Underhållsarbete hade utförts på merparten av de elva kulturarvsplatser vi
besökte, och några stödmottagare förklarade att fler arbeten hade planerats för
framtiden. I tre fall hade det varit nödvändigt att totalrenovera platsen på grund av
bristande underhåll i det förgångna. Detta visar på betydelsen av regelbundet
underhåll.
Förebyggande underhåll är också av grundläggande betydelse för att hantera
olika bevaranderisker som kulturplatser löper. Resultaten av vår enkät visar att
kulturarvsplatser är de platser som utsätts för de mest direkta hoten när det gäller
deras fysiska bevarande (se figur 4). De huvudsakliga risker som identifierades var
lokala förhållanden som påverkar platsens fysiska konstruktion (t.ex. regn, vind och
damm) och föroreningar. Men de största riskerna för stödmottagare, vilket gäller för
såväl ny kulturell infrastruktur som kulturarvsplatser, är faktorer som rör förvaltning
och institutionella frågor (t.ex. otillräckliga ekonomiska resurser och personalresurser
och avsaknad av en förvaltningsplan).
Figur 4 – Risker avseende bevarandet av kulturplatsen identifierade av
de 27 stödmottagarna i vårt urval (antal stödmottagare som identifierat
Förvaltning och institutionella faktorer
Lokala förhållanden som påverkar den fysiska
konstruktionen
Föroreningar
Plötsliga ekologiska eller geologiska händelser
Effekter av turism/besökare/rekreation
Klimatförändring och allvarliga väderfenomen
Annan mänsklig verksamhet
Byggnad och utveckling
Transportinfrastruktur
Sociala och kulturella användningsområden för kulturarv
Inga risker identifierade
Kulturarvsplats
Ny kulturell infrastruktur
Källa: Revisionsrätten, baserat på enkäten.
Underhåll och riskbedömning är inte finansieringskrav för de granskade Eruf-projekten
Ingen av de granskade stödmottagarna var tvungen att i samband med ansökan
om Eruf-finansiering visa hur deras plats skulle bevaras efter projektets slutförande
eller presentera en underhållsplan. Inte heller när det gällde kulturarvsplatser specifikt
ansågs frågan om hur brådskande de fysiska arbetena på platsen var som en viktig
faktor i Eruf-finansieringen, och i endast fyra urvalsförfaranden gynnades platser i
behov av mer brådskande arbete. Myndigheterna i medlemsstaterna krävde dock att
stödmottagarna skulle följa kvalitetsstandarder som fastställts i den nationella
lagstiftningen för de arbeten som skulle utföras under projektgenomförandet i 13 av
de 21 granskade urvalsförfarandena (se bilaga VI).
Enligt Eruf-förordningen ska det finnas nationella eller regionala riskbedömningar
för katastrofhantering som beaktar anpassning till klimatförändringar. Detta som en
förutsättning för att Eruf-medel från det tematiska målet att främja anpassning,
riskförebyggande och riskhantering i samband med klimatförändringar ska användas
ändamålsenligt och sparsamt. Eruf-ramen kräver inte att medlemsstaterna ska ta med
kulturarvsplatser, det vill säga de kulturplatser som är mer utsatta för naturliga faror, i
sina nationella eller regionala riskbedömningar. I en studie som kommissionen
genomförde nyligen angavs att skyddet av kulturarvet mot naturkatastrofer och
katastrofer orsakade av människan fortfarande påverkas negativt av det faktum att
kulturarvet ännu inte fullt ut ses, eller tas med, som en riskhanteringsprioritering i
nödsituationer 47. Tillsammans med medlemsstaterna angrep kommissionen detta
problem i december 2019 genom att utarbeta riktlinjer för rapportering om
katastrofriskhantering som bland annat hänvisar till kulturarvsplatser och som
uppmuntrar medlemsstaterna att rapportera, kartlägga och informera om de
potentiella konsekvenserna av katastrofrisker för kulturarvet 48. Det återstår att se hur
riktlinjerna kommer att tillämpas av medlemsstaterna.
En avvägning mellan hållbar turism och kulturarvsplatsers ekonomiska och sociala mål
Det är framför allt genom strategier för turismfrämjande som medlemsstaterna
skapar en socioekonomisk effekt med Eruf-investeringarna i kulturplatser (se
punkt 56). Effekterna av investeringarna mäts genom ”ökningen av antalet besökare
på platserna” (se punkt 66). Strategierna kan vara kontraproduktiva för bevarandet av
kulturarvsplatser som redan har problem med massturism. Att kulturarvsplatser
förstörs på grund av massturism var en risk som identifierades av 38 % av de förvaltare
av kulturarvsplatser som besvarade vår enkät (se figur 4). Vissa av de besökta
projekten har redan vidtagit åtgärder för att begränsa antalet turister eller för att
hantera turistströmmar på ett mer hållbart sätt (se ruta 7).
Europeiska kommissionen, Safeguarding Cultural Heritage from Natural and Man-Made
Disasters, A comparative analysis of risk management in the EU, 2018.
Riktlinjerna för rapportering antogs av kollegiet och offentliggjordes i december 2019
(EUT C 428, 20.12.2019, s. 8).
Ruta 7
Exempel på åtgärder som vidtagits för att kontrollera följderna av
överturism
Joanine-biblioteket från tidigt 1700-tal är en av juvelerna vid universitetet i
Coimbra i Portugal, som är ett av världens äldsta universitet och finns med på
Unescos världsarvslista. Det utformades arkitektoniskt så att en konstant
temperatur och luftfuktighet upprätthålls som gör att de litterära verken kan
bevaras. Eftersom turistbesök förekommer dagligen och den väldiga
huvudentrédörren i teak öppnas med jämna mellanrum uppstår ständiga
variationer i innetemperaturen och halten av damm, vilket påverkar det
långsiktiga bevarandet av de gamla, och ofta sällsynta, litterära verk som
biblioteket innehåller.
För att minska turistbesökens effekter har universitetet i Coimbra bytt
huvudingång till biblioteket. Tillträdet har också begränsats till grupper på högst
personer, som släpps in i omgångar på 20 minuter, och som får tillbringa högst
minuter i huvudsalen. Nyligen skaffade universitet även en anoxikammare som
återställer luftfuktighetsnivåer och avlägsnar svampar och parasiter från böcker
utan kemikalier.
Joanine-biblioteket i Coimbra i Portugal
© Fotograf: Henrique Patricio.
Arkitekt: Gaspar Ferreira.
Källa: Universitetet i Coimbra.
I liknande fall bör bevarandet av platsen prioriteras, oavsett vilken omedelbar
ekonomisk och social effekt det får. Men om insatserna på en plats inte förväntas få
sådana effekter, och även om de brådskar, kan Eruf för närvarande inte finansiera dem
(se punkterna 56–61). Det kan inte heller programmet Kreativa Europa. Detta var
tidigare möjligt genom Rafael-programmet 49 som löpte från 1997 till 2000 och bland
annat hade som mål att bevara, skydda och utveckla det europeiska kulturarvet.
EU har nyligen ökat sina ansträngningar för att säkerställa att kulturarvet bevaras
I efterdyningarna av branden i Notre-Dame-katedralen i Paris 2019 efterlyste de
kulturministrarna i EU:s medlemsstater att ett europeiskt nätverk för skydd av det
europeiska kulturarvet skulle inrättas och beslutade att skyddsfrågor ska ingå i EU:s
politik50.
Kommissionen tar indirekt upp riskreducering för kulturarvsplatser genom
förordningar om miljö- och energiprestanda. Medlemsstaterna har sedan 2012 varit
skyldiga att bedöma påverkan på kulturarvsplatser av offentliga och privata projekt
med betydande inverkan på miljön 51. Sedan 2018 ska medlemsstaterna ”[a]vseende
byggnader som genomgår större renoveringar  ta hänsyn till frågor som rör
brandsäkerhet och risker i samband med intensiv seismisk aktivitet” 52.
Inom ramen för Europaåret för kulturarv inledde kommissionen ett initiativ för
hotade kulturarv och gjorde en jämförande analys av riskhanteringspraxis i EU i syfte
att dela erfarenheter och främja samarbete mellan medlemsstater för att hantera
effekterna av naturkatastrofer eller katastrofer orsakade av människan på kulturarvet
(se punkt 73). Inom ramen för Europaåret för kulturarv har också en expertgrupp
under ledning av ICOMOS tagit fram kvalitetsprinciper för EU-finansierade projekt med
potentiell påverkan på kulturarvet 53. Kommissionen har ännu inte tagit ställning till om
och i så fall hur dessa principer ska beaktas på EU-nivå.
Beslut nr 2228/97/EG om att inrätta ett gemensamt åtgärdsprogram på kulturarvsområdet
(EGT L 305, 8.11.97, s. 31).
Se punkt 59.
Artikel 3 d i direktiv 2011/92/EU om bedömning av inverkan på miljön av vissa offentliga
och privata projekt, ändrat genom direktiv 2014/52/EU (EUT L 124, 25.4.2014, s. 1).
Artikel 7 i direktiv 2012/27/EG om energieffektivitet, ändrat genom direktiv (EU) 2018/844
(EUT L 156, 19.6.2018, s. 75).
ICOMOS, European Quality Principles for EU-funded interventions with potential impact
upon cultural heritage, 2019.
De granskade kulturplatserna är i allmänhet beroende av offentliga subventioner och
har få incitament att öka inkomsterna
De granskade kulturplatserna är i allmänhet beroende av offentliga subventioner
Vi analyserade självfinansieringsgraden för de kulturplatser där Eruf-projekten
hade slutförts. Självfinansieringsgraden är andelen driftskostnader som täcks av de
inkomster som platsens operativa verksamhet genererar (”egna medel”). Vi betraktar
en plats som finansiellt självförsörjande om de egna medlen överstiger eller är lika
med driftskostnaderna. Vi baserade vår bedömning på platsernas finansiella
räkenskaper från 2018.
Med undantag av tre projekt var ingen av de 21 granskade kulturplatser för vilka
uppgifter fanns tillgängliga finansiellt självförsörjande 2018. Kulturplatser är
huvudsakligen beroende av offentliga subventioner för sin drift. Privata donationer
förekommer men är av marginell betydelse. Vid åtta av de elva kulturplatser som fick
donationer 2018 täckte donationerna mindre än 3 % av respektive plats totala årliga
driftskostnader.
Kulturplatser är också starkt beroende av subventioner för att kunna finansiera
sina investeringskostnader. I 13 av de 23 granskade, slutförda projekten hade Erufinvesteringsprojekten finansierats helt med offentliga medel (från EU eller
nationella/lokala offentliga organ). Endast två av de granskade projekten fick privata
donationer. Beroendet av offentliga subventioner innebär en risk när det gäller den
kontinuerliga driften av kulturplatserna, eftersom de offentliga myndigheterna kan
minska finansieringen (se ruta 8).
Ruta 8
Exempel på risker för kulturplatser som är beroende av offentliga
subventioner och behovet av att diversifiera inkomstkällorna
Europeiska solidaritetscentrumet i Gdańsk i Polen har varit starkt beroende av
offentliga subventioner sedan det inrättades 2012. År 2019 minskade det polska
ministeriet för kultur och nationellt kulturarv sitt bidrag till kulturplatsen.
Solidaritetscentrumet var tvunget att genomföra gräsrotsfinansieringskampanjer
på sociala medier för att förbli finansiellt hållbart och för att kunna fortsätta att
bedriva sin normala verksamhet. Enligt centrumet hotas inte dess existens av det
ändrade offentliga stödet, men det har nödvändiggjort betydande ändringar av
verksamheten.
Den nuvarande finansieringsramen ger inte tillräckliga incitament till
inkomstgenerering
Enligt förordningen om gemensamma bestämmelser för 2014–2020 ska
stödmottagare ha den ekonomiska förmågan att genomföra det finansierade
projektet 54. I fråga om projekt som genererar nettoinkomster kräver förordningen om
gemensamma bestämmelser även att stödmottagarna i förväg ska uppskatta den
ström av inkomster och kostnader som genereras av EU-projektet för att identifiera
den eventuella del av investeringskostnaderna som behöver finansieras med EUmedel 55. Enligt förslaget till förordning om gemensamma bestämmelser för 2021–2027
måste medlemsstaterna kontrollera att stödmottagarna har de medel som krävs för att
täcka drifts- och underhållskostnaderna 56.
Projekts finansiella hållbarhet är därför ett kriterium som ofta används av
förvaltande myndigheter: det var ett krav i 20 av de 21 urvalsförfaranden som vi
granskade, antingen för att projekt skulle vara potentiellt berättigade till EU-stöd över
huvud taget (dvs. som ett tillåtlighetskriterium) eller för tilldelning av poäng när
projekt valdes ut (dvs. som ett urvalskriterium) – se bilaga V.
De förvaltande myndigheterna ansåg att de besökta projekten var finansiellt
hållbara eftersom det fanns en institutionell stödram som i princip garanterade deras
finansiella hållbarhet. Men i det stora flertalet fall var de faktiska
självfinansieringsgraderna lägre än vad som ursprungligen förutsågs i projektansökan
(se figur 5). Tre år efter projektslutförandet hade endast två av de 16 granskade
Artikel 125.3 d i förordningen om gemensamma bestämmelser.
Artikel 61 i förordningen om gemensamma bestämmelser.
Artikel 67.3 d i COM(2018) 375 final.
kulturplatser som det fanns uppgifter om uppnått resultatet enligt de ursprungliga
beräkningarna, medan självfinansieringsgraden för sex kulturplatser hade minskat med
över hälften. Detta förklaras av olika faktorer, till exempel överoptimistiska finansiella
prognoser eller stora förändringar av den ekonomiska modell som man planerat att
använda för kulturplatsen.
Figur 5 – Skillnader
mellan
självfinansieringsgrader
faktiska
och
%
%
Kulturplats nr 1
%
Kulturplats nr 2
%
Kulturplats nr 3
%
%
%
%
Kulturplats nr 8
%
%
Kulturplats nr 9
%
Kulturplats nr 10
Kulturplats nr 11
%
%
Kulturplats nr 13
%
Kulturplats nr 14
7%
2%
4%
%
%
%
%
%
%
Kulturplats nr 12
Kulturplats nr 16
%
6%
Kulturplats nr 7
Kulturplats nr 15
%
%
Kulturplats nr 5
%
%
%
Kulturplats nr 4
Kulturplats nr 6
prognostiserade
%
%
Faktisk självfinansieringsgrad (tre
år efter slutförandet eller, om
den tiden inte hade förflutit,
2018)
Förväntad självfinansieringsgrad
(tre år efter slutförandet)
Anm.: Diagrammet avser de slutförda projekt som det fanns uppgifter om. Den faktiska
självfinansieringsgraden hänför sig till tre år efter slutförandet av projektet eller, om den tiden inte hade
förflutit, till 2018.
Källa: Revisionsrätten, på grundval av stödmottagarnas finansiella räkenskaper.
44 
Eruf‐ramen ger inte stödmottagarna incitament att öka sina inkomster. Eruf‐
kraven på inkomstgenererande projekt innebär att ju högre nettoinkomster som 
projektet genererar, desto mindre blir EU‐stödet57. Men vid fyra besökta 
kulturarvsplatser var den ström av inkomster och kostnader som hade beräknats i 
förväg av begränsad relevans. Det berodde på att EU:s investeringar var inriktade på 
specifika delar av kulturplatsen (t.ex. på ett yttertak eller ett visst rum) som en del av 
platsens totala kostnader och intäkter måste tillskrivas, och den fördelningen 
baserades på uppskattningar och antaganden som inte alltid var tydliga. 
De urvalsförfaranden som vi granskade gav dessutom sällan incitament till 
inkomstgenererande verksamhet. Endast i ett fall kunde de sökande få upp till tre 
poäng om deras projekt ökade den aktuella andelen finansiering från privata källor. 
Alla intervjuade nationella experter angav att kulturplatserna inte utnyttjade 
inkomstgenererande verksamheters fulla potential, till exempel genom att starta 
souvenirbutiker, hyra ut lokaler eller utveckla strategier för biljettförsäljning eller ökad 
sponsorverksamhet (se tabell 4). 
Tabell 4 – Inkomstgenererande verksamheter som bedrevs av de besökta 
kulturplatserna i vårt urval, vilkas Eruf‐projekt hade slutförts vid 
tidpunkten för revisionen 
Biljett‐
försäljning 
(t.ex. besök, 
före‐
ställningar 
och ut‐
ställningar) 
Butiker 
(t.ex. 
souvenirer 
och 
böcker) 
Servering 
(t.ex. 
kafeteria och 
restaurang) 
Lokal‐
uthyr‐
ning 
Bidrags‐
kampanjer 
(t.ex. sponsring 
och donationer) 
OLIVA kreativfabrik 
X 
X 
X 
X 
 
Viana do Castelos 
kulturcenter 
X 
 
 
 
 
Katedralsleden 
X 
X 
 
 
X 
Pompeji 
X 
X 
X 
X 
X 
Villa Campolieto 
X 
 
 
X 
X 
San Carlo‐teatern 
X 
X 
X 
X 
X 
Sant Antonio‐
klostret 
 
 
 
 
 
Italien 
Portugal 
Medlemsstat/Projekt 
                                                       
  Se även punkt 97 i revisionsrättens särskilda rapport 06/2018. 
 
45 
Biljett‐
försäljning 
(t.ex. besök, 
före‐
ställningar 
och ut‐
ställningar) 
Butiker 
(t.ex. 
souvenirer 
och 
böcker) 
Servering 
(t.ex. 
kafeteria och 
restaurang) 
Lokal‐
uthyr‐
ning 
Bidrags‐
kampanjer 
(t.ex. sponsring 
och donationer) 
Polens nationella 
radiosymfoni‐
orkester 
X 
 
 
X 
 
Solidaritets‐
centrumet 
X 
X 
X 
X 
X 
Paviljongen Fyra 
kupoler 
X 
X 
 
X 
X 
Polen 
Medlemsstat/Projekt 
Källa: Revisionsrätten. 
 
 
 
På projektnivå var de granskade kulturplatsernas förmåga och incitament att
diversifiera sina egna medel ännu i många fall rättsligt och finansiellt begränsade.
Enligt de experter vi intervjuade får kulturplatser ofta motstridiga incitament. Till
exempel kan generering av ytterligare inkomster leda till efterföljande nedskärningar
av den offentliga finansieringen. I genomsnitt har kulturplatser som är administrativt
och finansiellt självständiga högre självfinansieringsgrad (se figur 6).
Figur 6 – Faktisk självfinansieringsgrad hos slutförda, granskade projekt
Självständiga platser
Icke självständiga platser
%
%
Anm.: Diagrammet avser de slutförda projekt som det fanns uppgifter om. Den faktiska
självfinansieringsgraden hänför sig till tre år efter slutförandet av projektet eller, om den tiden inte hade
förflutit, till 2018.
Källa: Revisionsrätten, på grundval av stödmottagarnas finansiella räkenskaper.
En avvägning mellan finansiell hållbarhet och uppnåendet av kulturella och sociala mål
Finansiella begränsningar gör att man måste välja. Valen kan leda till lägre
investeringar i bevarandet av den fysiska infrastrukturen, till ett minskat utbud av
kulturverksamheter eller till begränsningar av tillträdet till kulturplatsen på grund av
att man har behövt höja inträdesavgifterna. Det gäller att hitta en balans mellan vad
som förväntas av kulturplatser socialt och kulturellt och vad de faktiskt kan
åstadkomma (se ruta 9).
Ruta 9
Att kombinera tillgång till kultur och finansiell stabilitet
Museet Louvre-Lens erbjöd fritt inträde till sin permanenta utställning
(”Tidsgalleriet”) och till en av sina tillfälliga utställningshallar (”Glaspaviljongen”)
för att öka tillgången till kultur och locka nya besökare. Enligt museet ökade denna
åtgärd det totala antalet besökare 58 (14 % av besökarna skulle inte ha besökt
museet om de hade varit tvungna att betala en inträdesavgift) men begränsade
dess finansiella självständighet genom att självfinansieringsgraden minskades 59
(18 % i stället för förväntade 27 %). Gratis inträde har hittills kunnat behållas tack
vare att de lokala myndigheterna åtagit sig att täcka museets driftsunderskott.
När projekten har slutförts är medlemsstaternas projektövervakning begränsad
Enligt den rättsliga grunden60 ska stödmottagarna upprätthålla EU-projektets
karaktär och mål under en varaktighetsperiod på fem år. Överträdelser av dessa
skyldigheter kan leda till finansiella korrigeringar och återvinningar av de beviljade EUmedlen. EU:s rättsliga ram anger inte hur de förvaltande myndigheterna i
medlemsstaterna ska säkerställa efterlevnad av dessa krav. Det är medlemsstaternas
ansvar att fastställa adekvata övervakningsarrangemang.
De förvaltande myndigheterna övervakar projekten i första hand under
genomförandefasen. Trots att målvärdena för omkring en fjärdedel av de
resultatindikatorer som fastställts för de slutförda projekten i vårt urval inte hade
uppnåtts vid slutförandet (se även figur 3) fick det inga finansiella konsekvenser för
stödmottagarna. Vi har i en tidigare rapport angett att incitamentsmekanismerna ska
tillämpas och leda till verkliga ekonomiska fördelar eller sanktioner 61. ICOMOS har
angett att de övervakningsförfaranden som fastställts av EU och medlemsstaterna för
EU-finansierade projekt inte tar tillräcklig hänsyn till kultursektorns särdrag och lägger
för stor vikt vid finansiella aspekter utan en ordentlig bedömning av projektens faktiska
kvalitet och kulturella påverkan (se ruta 10).
Louvre Lens, 5 ans de gratuité de la galerie du temps et du pavilion de verre: bilan et
perspectives, mars 2018, s. 12.
Franska regionala revisionsorganet i Nord–Pas-de-Calais/Picardie, Établissement public de
coopération culturelle « Louvre-Lens » Exercices 2011 et suivants, Relevé d’observations
définitives, 2015, s. 9.
Artikel 71 i förordningen om gemensamma bestämmelser.
Punkterna 54–56 i revisionsrättens briefingdokument om en prestationsinriktad
sammanhållningspolitik, juni 2019.
Ruta 10
Exempel på bristande fokus på kulturella aspekter
Världsarvet i Pompeji beviljades Eruf-medel på cirka 78 miljoner euro till skydd
och främjande. Arbeten utfördes på olika ställen på platsen. För vårt
revisionsbesök valde vi ut Efebo-huset, som slutfördes i december 2015.
Bland annat restaurerades husets ”sommar-triclinium”, en romersk matsal som
användes sommartid med utsikt över trädgården under en pergola som bärs upp
av fyra kolonner. Den förvaltande myndigheten besökte Efebo-huset för att
verifiera de redovisade kostnaderna. Myndighetens rapport bekräftade att
arbetena hade slutförts.
Tre år efter arbetenas slutförande hade byggnaden skador på ett antal ställen.
Under en övervakningskontroll som stödmottagaren gjorde drog experter
slutsatsen att byggnaden hade underminerats av det mycket stora antalet
besökare som hade tillträde till triclinium och av avsaknaden av skydd på
byggnadens samtliga sidor. Ett skydd av polykarbonat hade finansierats av det
granskade Eruf-projektet men det hade förvarats i ett magasin och aldrig
monterats. Det monterades i början av 2019 i samband med underhållsarbeten,
tre år efter det att projektet hade slutförts. Detta fel skadade sommar-tricliniums
fysiska infrastruktur.
Sommar-triclinium, 1927
Källa: Scheda ispettiva, Casa dell’Efebo I 7, 11, från Parco Archeologico di Pompei.
Sommar-triclinium, januari 2016, efter slutförandet av det granskade Erufprojektet 2015
Källa: Relazione tecnica, Casa dell’Efebo, januari 2016, från Parco Archeologico di Pompei.
Sommar-triclinium, april 2019, under revisionsbesöket
Källa: Revisionsrätten.
Efter projektens slutförande säkerställer inte övervakningssystemen i de besökta
medlemsstaterna att projektens prestation kontrolleras regelbundet. Under den
femåriga varaktighetsperioden kan prestationen kontrolleras på ad hoc-basis, efter
nationellt gottfinnande. Därefter övervakas inte projektens prestation.
På projektnivå hade endast en av de besökta kulturplatserna genomgått en
efterhandsbedömning för analys av Eruf-projektets ekonomiska, sociala eller kulturella
effekter.
Vad beträffar kulturarvsplatser står Erufs övervakningsarrangemang i tydlig
kontrast till de arrangemang som införts för Unesco och Europarådets kulturvägar
samt av kommissionen själv när det gäller platser som fått Europeiska
kulturarvsmärket. Eruf tillhandahåller medel men kräver ändå inte att projekten ska
övervakas regelbundet efter det att de har slutförts. Medlemsstaternas praxis
härvidlag varierar kraftigt under den femåriga varaktighetsperioden. När det gäller
programperioden 2014–2020 övervakar två av de besökta medlemsstaterna vissa
projekt på plats, medan en medlemsstat endast gör administrativa kontroller på
grundval av rapporter som stödmottagarna lämnar in. I motsats till det krävs enligt de
tidigare nämnda internationella utmärkelserna att övervakning ska utföras
systematiskt, trots att de inte nödvändigtvis tillhandahåller medel (se bilaga VII).
Slutsatser och rekommendationer
Den samlade slutsatsen av revisionen är att det saknas en lämplig ram som
garanterar att Eruf-investeringar i kulturplatser blir ändamålsenliga och hållbara.
Bristande fokus och begränsad samordning när det gäller EU:s
investeringar i kulturplatser
Fördragen fastställer som överordnat mål att EU ska respektera rikedomen hos
sin kulturella mångfald och sörja för att det europeiska kulturarvet skyddas och
utvecklas. Kultur är huvudsakligen medlemsstaternas behörighet. Unionen kan endast
uppmuntra till samarbete mellan medlemsstater och stödja eller komplettera deras
insatser (punkterna 05–16).
Kultur behandlas inte i kommissionens övergripande Europa 2020-strategi. EU:s
grundläggande strategiska ram för kultur består av gemensamma strategiska mål som
vägleder EU:s insatser på kulturområdet. Målen fastställs i kommissionens agendor för
kultur och preciseras i rådets arbetsplaner för kultur. Denna ram är komplex. Den
förekommer parallellt med många olika allmänna strategiska EU-ramar och EU-mål
med överlappande perioder och flera ansvarsnivåer. De strategiska mål som
kommissionen har fastställt omvandlas inte till tydliga operativa mål, och det finns inga
bestämmelser om övervakning av måluppfyllelse eller indikatorer för att mäta
framsteg. Enligt kommissionen är det fortfarande en utmaning att omvandla mål till
politiska beslut på medlemsstatsnivå (punkterna 17–22).
Den strategiska ramen för kultur återspeglas dessutom endast delvis i EU:s
finansiering. Kulturella aspekter införlivas, eller ”integreras”, i olika politikområden och
betraktas framför allt som en resurs som bidrar till uppnåendet av andra EUprioriteringar och EU-mål genom olika EU-fonder. Men av de tolv EU-fonder som
potentiellt skulle kunna stödja kultur som vi analyserade hänvisar endast förordningen
om Kreativa Europa, som är en liten fond sett till budgeten, till kommissionens agenda
från 2007. Det här gör att nyttan med agendan kan ifrågasättas (punkterna 23–24).
Kommissionen har tagit åtskilliga initiativ för att främja kulturplatser, men EU:s
kulturinitiativ har mycket begränsad effekt på stödmottagares tillgång till Eruf-medel.
Eruf-förordningen fastställer högre finansieringsgränser för Unescos världsarvsplatser,
men det finns inga sådana bestämmelser för kulturplatser som har en EU-utmärkelse
eller som deltar i ett av EU:s kulturinitiativ. Samordningen mellan EU:s fonder för
investeringar i kulturplatser är också mycket begränsad (punkterna 25–36).
På EU-nivå finansieras infrastrukturinvesteringar framför allt genom Eruf. Eruf är
en viktig källa till finansiering av investeringar i kulturplatser för omkring en tredjedel
av medlemsstaterna. Men Eruf prioriterar inte investeringar i kulturplatser utan stöder
ett annat fördragsmål: främjandet av social och ekonomisk sammanhållning. Vi fann
exempel på att medlemsstater hade tagit initiativ till finansiering av kulturplatser och
utveckling av finansieringssystem som byggde på privata medel (punkterna 37–51).
Rekommendation 1 – Förbättra den nuvarande strategiska
ramen för kultur i enlighet med de befogenheter som anges i
fördragen
Kommissionen bör med beaktande av sina befogenheter föreslå att
medlemsstaterna ska fastställa tydliga strategiska och operativa mål i nästa
arbetsplan för kultur. Målen bör övervakas regelbundet genom indikatorer med
målvärden och delmål.
Ansvaret för genomförandet av målen bör fastställas och fördelas, bland annat
lämplig samordning inom kommissionen.
Kommissionen bör identifiera och ge intressenter exempel på god praxis för hur
EU-finansierade kulturprojekt ska utformas, väljas ut, finansieras, genomföras och
övervakas/följas upp. I detta skulle framför allt upprättande av underhållsplaner,
utveckling av sociala verksamheter och kulturplatsers deltagande i EU-initiativ
kunna ingå.
Tidsram: Senast i december 2022.
Rekommendation 2 – Uppmuntra användning av privata medel
för att skydda Europas kulturarv
För att bättre försöka uppfylla EU-fördragets mål att skydda det europeiska kulturarvet
bör kommissionen
samla god praxis när det gäller alternativa finansieringskällor i medlemsstaterna,
tillsammans med medlemsstaterna undersöka möjligheten att utveckla ett system
som bygger på privata källor till finansiering av kulturarvsplatser,
samordna sådana potentiella initiativ med andra EU-initiativ på kulturområdet
(t.ex. europeiska kulturarvsmärket och europeiska kulturhuvudstäder).
Tidsram: Senast i december 2022.
Varierande ändamålsenlighet och hållbarhet hos de granskade Erufprojekten
Trots EU:s ambition att öka kulturinsatsernas sociala effekter är målen för Erufs
operativa program och projekt mestadels ekonomiska. Investeringar i kulturplatser
betraktas som en resurs för att öka konkurrenskraften eller utveckla lokala områden.
Kulturella aspekter ägnades minst uppmärksamhet i de granskade operativa
programmen, även i de fall då de tydligt angavs som mål. De förvaltande
myndigheterna inom Eruf ansåg ofta att kulturella aspekter inte var relevanta när de
valde ut projekt (punkterna 52–61).
Projektens prestation kunde inte bedömas för alla granskade projekt som hade
slutförts. Projekten var operativa vid tidpunkten för revisionen, men vi fann flera
brister i urvalet och rapporteringen av indikatorer som begränsar möjligheten att
använda de rapporterade uppgifterna för att dra slutsatser om projektens prestation.
På grund av karaktären på Erufs resultatindikatorer är dessutom uppfyllelsen av de
operativa programmens mål inte alltid direkt beroende av enskilda projekts prestation
(punkterna 62–67).
Eruf-kraven gäller inte det fysiska bevarandet av kulturplatser som fått
finansiering. Trots kulturarvsplatsers fortlöpande behov av underhåll och de många
bevaranderisker som de löper, behövde inget av de granskade Eruf-projekten visa hur
kulturplatsen skulle bevaras efter projektets slutförande eller presentera en
underhållsplan i samband med ansökan om EU-medel. Vidare kan varken Eruf eller
Kreativa Europa finansiera bevarandet av utsatta kulturplatser om inte arbetet
förväntas ha direkta ekonomiska och sociala effekter. Detta var tidigare möjligt genom
Rafael-programmet. För platser som redan har problem med massturism kan
skapandet av ekonomiska effekter, ofta genom strategier för turismfrämjande, vara
kontraproduktivt för bevarandet av dem (punkterna 68–75).
EU har nyligen ökat sina ansträngningar för att säkerställa att kulturarvet
bevaras. Men på medlemsstatsnivå kräver inte Eruf-ramen att medlemsstaterna ska
integrera kulturarvsplatser, det vill säga de kulturplatser som är mest utsatta när det
gäller naturkatastrofer, i de nationella eller regionala riskbedömningar som ska göras
enligt EU:s lagstiftning (punkterna 76–78).
De granskade kulturplatserna är i allmänhet beroende av offentliga
subventioner för sin drift och finansiering av investeringskostnader. Eruf-ramen ger
inte stödmottagarna incitament att öka sina inkomster. Eruf-kraven på
inkomstgenererande projekt innebär att ju högre nettoinkomster som projektet
genererar, desto mindre blir EU-stödet. De urvalsförfaranden som vi granskade gav
dessutom sällan incitament till inkomstgenererande verksamhet (punkterna 79–88).
När projekten har slutförts är projektövervakningen begränsad.
Övervakningssystemen i de besökta medlemsstaterna möjliggör kontroll av projektens
prestation på ad hoc-basis under den varaktighetsperiod på fem år som krävs enligt
EU:s lagstiftning, men därefter övervakas inte prestationen mer. I de granskade
projekten påverkade inte heller projektens prestation storleken på det Eruf-belopp
som stödmottagarna erhöll (punkterna 89–93).
Rekommendation 3 – Stärk den finansiella hållbarheten för
kulturplatser som finansieras av Eruf
För att inte avskräcka stödmottagare från att öka sina egna inkomster bör
kommissionen undersöka och föreslå förenklade former av stöd för Eruf-investeringar i
kulturplatser.
För att minska beroendet av offentliga subventioner bör Eruf-finansieringen under den
fas då projekten väljs ut gynna projekt som innehåller planer för att förbättra
kulturplatsers finansiella självförsörjning (t.ex. diversifiering av och ökad användning av
egna inkomstmedel).
Tidsram: I tid till förhandlingarna om de operativa programmen för programperioden
2021–2027.
Rekommendation 4 – Vidta mer specifika åtgärder för att
bevara kulturarvsplatser
När kommissionen förhandlar om operativa program bör den rekommendera
medlemsstaterna att inkludera kulturarvsplatser i de nationella eller regionala
riskhanteringsplaner för katastrofer som föreskrivs i den föreslagna förordningen om
gemensamma bestämmelser. Det skulle uppmuntra dem att identifiera de
bevaranderisker som kulturarvsplatser löper och planera lämpliga riskreducerande
åtgärder.
Tidsram: I tid till förhandlingarna om de operativa programmen för programperioden
2021–2027.
Denna rapport antogs av revisionsrättens avdelning II, med ledamoten Iliana Ivanova
som ordförande, vid dess sammanträde i Luxemburg den 26 februari 2020.
För revisionsrätten
Klaus-Heiner Lehne
ordförande
Bilagor
Bilaga I – Översikt över offentliga utgifter för kulturella tjänster
Utgifter för kulturella tjänster per invånare och som andel av de totala offentliga
utgifterna
euro
Lettland
3,0 %
Estland
2,6 %
Ungern
2,6 %
Malta
2,2 %
Litauen
2,0 %
Polen
1,7 %
Kroatien
1,6 %
Bulgarien
1,6 %
Slovenien
1,5 %
Tjeckien
1,5 %
Danmark
1,3 %
Luxemburg
1,2 %
Frankrike
1,2 %
Slovakien
1,1 %
Österrike
1,1 %
Spanien
1,1 %
Rumänien
1,0 %
Sverige
1,0 %
Belgien
1,0 %
Finland
1,0 %
Nederländerna
1,0 %
EU-28
1,0 %
Tyskland
0,9 %
Irland
0,8 %
Cypern
Belopp (i euro) per person i
befolkningen som gått till kulturella
tjänster
0,7 %
Förenade kungariket
0,6 %
Italien
0,6 %
Portugal
Grekland
0,5 %
0,3 %
Kulturella tjänsters andel av de totala
offentliga utgifterna
Kapitalinvesteringar i kulturella tjänster (absoluta belopp och som andel av de totala
offentliga utgifterna för kulturella tjänster)
miljoner euro
1 000
2 000
1 500
2 500
3 000
Luxemburg
%
Estland
%
Italien
%
Ungern
%
Malta
%
Lettland
%
Polen
%
Portugal
%
Frankrike
%
Cypern
%
Tjeckien
%
Litauen
%
Genomsnitt EU-28
%
Slovenien
%
Tyskland
%
Slovakien
%
Förenade…
%
Rumänien
%
Belgien
%
Irland
%
Österrike
%
Nederländerna
%
Danmark
%
Finland
9%
Spanien
9%
Bulgarien
7%
Kroatien
Grekland
Sverige
3 500
6%
Totala kapitalinvesteringar i kulturella
tjänster
Kapitalinvesteringarnas andel av de offentliga
utgifterna för kulturella tjänster
4%
3%
Anm.: Vi har använt Eurostats data om offentliga utgifter för kulturella tjänster (COFOG: GF08.2) för att
uppskatta medlemsstaternas investeringar i kulturplatser. Detta är den bästa uppskattning som finns
tillgänglig. Kapitalinvesteringar i kulturella tjänster inbegriper: investeringsbidrag (D92), fasta
bruttoinvesteringar (P.51g) och anskaffning minus avyttringar av icke finansiella icke producerade
tillgångar (NP). Siffrorna representerar de belopp som användes 2017 av nationella och lokala
myndigheter (offentliga utgifter).
Källa: Revisionsrätten, på grundval av Eurostat, General government expenditure by function (COFOG),
onlinedatakod: [gov_10a_exp].
Bilaga II – Översikt över EU-fonder med kulturella mål
Program
Programnamn
Ansvarigt GD
Antal
allmänna
mål
… där kultur Antal särskilda mål eller
nämns
investeringsprioriteringar
… med
kulturellt
innehåll
Hänvisar
Medel
till EU:s
tillgängliga för
agenda
investeringar i
för
kulturplatser?
kultur?
Rubrik 1a i den fleråriga budgetramen: Konkurrenskraft för tillväxt och sysselsättning
Horisont 2020
FSE
Erasmus+
Efsi
Ramprogrammet för
GD Forskning och
forskning och
innovation
innovation
Fonden för ett
GD Transport och
sammanlänkat Europa
rörlighet
EU:s program för allmän
GD Utbildning,
utbildning,
ungdom, idrott och
yrkesutbildning,
kultur
ungdom och idrott
Europeiska fonden för
strategiska
GD Ekonomi och
investeringar/EUfinans
garantin
Nej
Nej
Nej
Nej
Nej
Nej
Nej
Ja
Nej
Ja
Nej
Nej
Nej
Nej
Rubrik 1b i den fleråriga budgetramen: Ekonomisk, social och territoriell sammanhållning
GD Regional- och
stadspolitik
GD Sysselsättning,
ESF
Europeiska socialfonden socialpolitik och
inkludering
GD Regional- och
Sammanhållningsfonden Sammanhållningsfonden
stadspolitik
Eruf
Europeiska regionala
utvecklingsfonden
Program
Programnamn
Ansvarigt GD
Antal
allmänna
mål
… där kultur Antal särskilda mål eller
nämns
investeringsprioriteringar
… med
kulturellt
innehåll
Hänvisar
Medel
till EU:s
tillgängliga för
agenda
investeringar i
för
kulturplatser?
kultur?
Rubrik 2 i den fleråriga budgetramen: Hållbar tillväxt: naturresurser
Ejflu
EHFF
Life
Europeiska
jordbruksfonden för
landsbygdsutveckling
Europeiska havs- och
fiskerifonden
Program för miljö och
klimatpolitik
GD Jordbruk och
landsbygdsutveckling
Nej
Ja
GD Havsfrågor och
fiske
Nej
Ja
GD Miljö
Nej
Nej
Nej
Nej
Ja
Nej
Rubrik 3 i den fleråriga budgetramen: Säkerhet och medborgarskap
Ett Europa för
medborgarna
Kreativa Europa
Ett Europa för
medborgarna
Programmet Kreativa
Europa
GD Migration och
inrikes frågor
GD Utbildning,
ungdom, idrott och
kultur
Källa: Revisionsrätten, på grundval av EU-förordningar, relevanta inbjudningar att lämna förslag och 2007 års europeiska agenda för kultur som antogs genom rådets resolution av
den 16 november 2007.
Bilaga III – Lista över granskade insatsområden och tillhörande operativa program
Granskade operativa program
Programperiod
Medlemsstat
Titel
Granskade insatsområden (IO)
2014PT16M2OP002
Regionen Mellersta Portugal
IO 7. Bekräfta territoriernas
hållbarhet
IO 9. Stärka det urbana nätverket
Italien
2014IT16RFOP001
Kultur och utveckling
IO 1. Öka kulturanslagen
Polen
2014PL16M1OP001
Infrastruktur och miljö
IO VIII. Skydd av kulturarvet och
utveckling av kulturresurser
Frankrike
2014FR16M0OP012
Nord-Pas-de-Calais
IO 4. Öka regionens kapacitet att
anpassa sig till förändringar och även
dess attraktivitet och synlighet
Kroatien
2014HR16M1OP001
Konkurrenskraft och
sammanhållning
IO 6. Miljöskydd och resursernas
hållbarhet
Rumänien
2014RO16RFOP002
Regionalt operativt program
IO 5. Förbättring av stadsmiljön och
bevarande, skydd och hållbart
nyttjande av kulturarvet
Tyskland
2014DE16RFOP008
Mecklenburg-Vorpommern
IO 4. Främja integrerad och hållbar
stadsutveckling
Portugal
2014–2020
Operativt program
Programperiod
Medlemsstat
Titel
Granskade insatsområden (IO)
2007PT161PO002
Regionen Norra Portugal
IO II. Ekonomiskt främjande av
specifika resurser
IO III. Stärka den regionala
dimensionen
IO IV. Lokal och urban
sammanhållning
Italien
2007IT161PO001
Kultur-, natur- och
turistattraktioner
IO 1. Främjande och integrering av
kultur- och naturarvet på regional
nivå
Polen
2007PL161PO002
Infrastruktur och miljö
IO XI. Kultur och kulturarv
Frankrike
2007FR162PO017
Nord-Pas-de-Calais
IO 4. Territoriell dimension
Portugal
2007–2013
Operativt program
Kroatien
2007HR161PO003
Regional konkurrenskraft
IO 1. Utveckling och uppgradering av
den regionala infrastrukturen och
ökning av regionernas
attraktionskraft
IO 2. Stärkande av den kroatiska
ekonomins konkurrenskraft
Rumänien
2007RO161PO001
Regionalt operativt program
IO 5. Hållbar utveckling och hållbart
främjande av turism
Tyskland
2007DE162PO010
Niedersachsens regionala program
(utom Lüneburg)
IO 3. Stöd till den särskilda
infrastrukturen för hållbar tillväxt
Bilaga IV – Lista över granskade projekt
Medlems
-stat
Projektnamn
Programperiod
Besökt
Ja/Nej
Typ av plats
Grad av
självständighet
Läget vid
tidpunkten
för
revisionen
Totalt Erufbelopp (mn
EUR)*
Antal
outputindikatorer
Antal
resultatindikatorer
Portugal
Coimbras
universitet
2014–2020
Ja
Kulturarvsplats
Självständigt
Pågår
e.t.
Portugal
Convento
Abrantes
2014–2020
Ja
Kulturarvsplats
Ej självständigt
Pågår
e.t.
Portugal
OLIVA
2007–2013
Ja
Ny kulturell
infrastruktur
Ej självständigt
Slutfört
6,9
Portugal
Rota das
Catedrais
2007–2013
Ja
Kulturarvsplats
Självständigt
Slutfört
1,9
Portugal
Centro Cultural
de Viana
2007–2013
Ja
Ny kulturell
infrastruktur
Ej självständigt
Slutfört
10,7
Polen
Jasna Góra
Częstochowa
2014–2020
Ja
Kulturarvsplats
Självständigt
Slutfört
4,1
Polen
Toruń – gamla
staden
2014–2020
Ja
Kulturarvsplats
Ej självständigt
Pågår
e.t.
Medlems
-stat
Typ av plats
Grad av
självständighet
Läget vid
tidpunkten
för
revisionen
Totalt Erufbelopp (mn
EUR)*
Antal
outputindikatorer
Antal
resultatindikatorer
Projektnamn
Programperiod
Besökt
Ja/Nej
Polen
Europeiska
solidaritetscentr
umet i Gdańsk
2007–2013
Ja
Ny kulturell
infrastruktur
Självständigt
Slutfört
24,9
Polen
Paviljongen Fyra
kupoler
Wrocław
2007–2013
Ja
Kulturarvsplats
Självständigt
Slutfört
12,2
Polen
NOSPR Katowice
2007–2013
Ja
Ny kulturell
infrastruktur
Självständigt
Slutfört
33,7
Italien
Palazzo
Lanfranchi,
Matera
2014–2020
Ja
Kulturarvsplats
Ej självständigt
Pågår
e.t.
Italien
Ex Convento di
Sant’Antonio
2014–2020
Ja
Kulturarvsplats
Ej självständigt
Slutfört
2,7
Italien
Teatro di San
Carlo di Napoli
2007–2013
Ja
Kulturarvsplats
Självständigt
Slutfört
19,7
Italien
Villa Campolieto
2007–2013
Ja
Kulturarvsplats
Självständigt
Slutfört
4,2
Medlems
-stat
Projektnamn
Programperiod
Besökt
Ja/Nej
Typ av plats
Grad av
självständighet
Läget vid
tidpunkten
för
revisionen
Totalt Erufbelopp (mn
EUR)*
Antal
outputindikatorer
Antal
resultatindikatorer
Italien
Pompeji (Casa
dell’Efebo)
2007–2013
Ja
Kulturarvsplats
Självständigt
Slutfört
0,6
Rumänien
Mănăstirea
Moldovita
2007–2013
Nej
Kulturarvsplats
Självständigt
Slutfört
1,1
Rumänien
Muzeul
Judetean Buzău
2007–2013
Nej
Kulturarvsplats
Självständigt
Slutfört
4,7
Rumänien
Palatul
Patriarhiei,
Bukarest
2007–2013
Nej
Kulturarvsplats
Självständigt
Slutfört
12,6
Frankrike
Centre
Eurorégional
des cultures
urbaines (Lille)
2007–2013
Nej
Ny kulturell
infrastruktur
Ej självständigt
Slutfört
3,6
Frankrike
Halle au sucre
(Dunkerque)
2007–2013
Nej
Ny kulturell
infrastruktur
Ej självständigt
Slutfört
6,9
Frankrike
Musée du
Louvre Lens
2007–2013
Nej
Ny kulturell
infrastruktur
Självständigt
Slutfört
35,0
Medlems
-stat
Projektnamn
Programperiod
Besökt
Ja/Nej
Typ av plats
Grad av
självständighet
Läget vid
tidpunkten
för
revisionen
Totalt Erufbelopp (mn
EUR)*
Antal
outputindikatorer
Antal
resultatindikatorer
Kroatien
Muzej Rijeka
(Karlovac)
2007–2013
Nej
Ny kulturell
infrastruktur
Självständigt
Slutfört
4,7
Kroatien
Kneževe palače
(Zadar)
2007–2013
Nej
Kulturarvsplats
Ej självständigt
Slutfört
4,7
Kroatien
Ivanina kuća
bajke (Ogulin)
2007–2013
Nej
Ny kulturell
infrastruktur
Självständigt
Slutfört
0,9
Tyskland
Dom-Museum
Hildesheim
2007–2013
Nej
Kulturarvsplats
Ej självständigt
Slutfört
3,5
Tyskland
Kulturetage
Oldenburg
2007–2013
Nej
Ny kulturell
infrastruktur
Självständigt
Slutfört
2,0
Tyskland
Sprengel
Museum
Hannover
2007–2013
Nej
Ny kulturell
infrastruktur
Ej självständigt
Slutfört
11,6
Anm.: Indikatorerna avser projektens ekonomiska, sociala eller kulturella dimension.
Källa: Revisionsrätten.
Bilaga V – Översikt över de 21 granskade urvalsförfarandena
Tabellen ger en översikt över de krav som stödmottagarna enligt de förvaltande myndigheterna skulle uppfylla när de ansökte om Eruf-finansiering. I tabellen anges om
kraven betraktades som tillåtlighets- eller urvalskriterium. Tillåtlighetskriterierna inbegriper kriterier för stödberättigande och måste vara uppfyllda för att
stödmottagarna ska anses berättigade till finansiering. Uppfyllelse av ett urvalskriterium innebär en fördel för stödmottagaren (i form av extra poäng) men är inte
obligatoriskt.
Programperioden 2007–2013
Förvaltande myndigheters krav/Andel
urvalsförfaranden där stödmottagarna var skyldiga
att uppfylla kravet
Projektets ekonomiska effekt
Projektets sociala effekt
Ökning av antalet besökare
Införlivande i en lokal utvecklingsstrategi
Projektets kulturella effekt
- Projektets kulturella kvalitet
- Förekomst av ett kulturmärke (Unescos eller ett
nationellt märke)
- Deltagande i EU-initiativ (eller märken)
- Akut behov av fysiska åtgärder
- Effekt på anseendet och kulturarvsfrämjandet
Restaurering/Underhåll av platsen
- Kvalitet på de arbeten som ska utföras
- Fysiskt underhåll och underhållsplaner
Finansiell hållbarhet
- Rapportens kostnadseffektivitet
- Finansiell hållbarhet kan påvisas
Källa: Revisionsrätten.
Tillåtlighetskriterier
Urvalskriterier
Programperioden 2014–2020
Högsta
genomsnittliga
tilldelade viktning (i
förekommande fall)
%
%
%
%
Tillåtlighetskriterier
Urvalskriterier
Högsta
genomsnittliga
tilldelade viktning (i
förekommande fall)
%
%
%
%
e.t.
%
%
%
e.t.
%
e.t.
e.t.
%
8%
%
0%
%
e.t.
%
%
6%
7%
Ett krav i mellan 75 och 100 % av alla granskade urvalsförfaranden
Ett krav i mellan 50 och 75 % av alla granskade urvalsförfaranden
Ett krav i mellan 25 och 50 % av alla granskade urvalsförfaranden
Ett krav i mindre än 25 % av alla granskade urvalsförfaranden
Inte ett krav i något granskat urvalsförfarande
Bilaga VI – Lista över de viktigaste policydokumenten avseende
kulturplatser
Dokumentets titel
Typ av dokument
Datum
Behovet att framhäva kulturarvet i EU:s politik
Rådets slutsatser
Europeisk ram för åtgärder för kulturarv
Arbetsdokument från
kommissionens avdelningar
Europaåret för kulturarv
Europaparlamentets och
rådets beslut (EU) 2017/864
En enhetlig EU-politik för den kulturella och
kreativa sektorn
Parlamentets resolution
En integrerad kulturarvsstrategi för Europa
Parlamentets resolution
En integrerad kulturarvsstrategi för Europa
Meddelande från
kommissionen
Kartläggning av kulturarvsrelaterade åtgärder
i EU:s politikområden, program och
verksamheter
Meddelande från
kommissionen
Kulturarvet som en strategisk resurs för ett
hållbart Europa
Rådets slutsatser
Att främja de kulturella och kreativa
sektorerna för att främja tillväxt och
sysselsättning i EU
Meddelande från
kommissionen
Källa: Revisionsrätten.
Bilaga VII – Viktigaste kännetecken för europeiska
kulturarvsmärket, världsarvslistan och kulturvägar
EU:s europeiska
kulturarvsmärke1)
Unescos världsarv2)
Europarådets
kulturvägar3)
Medlemsstaterna
Konventionsstaterna
Europarådet, utökat
delavtal om kulturvägar
Antal platser/nätverk
med utmärkelser
platser
platser, varav 373 i
EU
inrättade europeiska
nätverk
Antal länder med
platser/nätverk med
utmärkelser
Skydda kulturarv med
enastående universellt
värde
Främja en gemensam
europeisk identitet och
gemensamma
europeiska värderingar,
interkulturell dialog, ett
europeiskt minne,
europeisk historia och
europeiskt kulturarv
Europeisk betydelse
Enastående universellt
värde
Europeiskt värde +
transnationell
dimension + europeiskt
minne, europeisk
historia och europeiskt
kulturarv
Övervakningsintervall
Vart fjärde år
Vart sjätte år
Vart tredje år
Utvärdering på platsen
Baserat på
självrapportering
Baserat på
självrapportering
Görs av en oberoende
expert
Inrättades
Ansvariga myndigheter
Främja europeisk
Viktigaste övergripande integration, historia och
principer
kultur samt europeiska
värden
Huvudkriterier för
tilldelning av
utmärkelsen
Aspekter som framför
allt övervakas
Feedback kring
Bevarandestatus,
utmärkelsen (fördelar,
förvaltning,
antal besökare etc.),
övervakningsförfaranden,
verksamheter till nästa verksamheter, risker, ny
period och
lagstiftning och effekter av
kommunikationsbehov
utmärkelsen
Teman, verksamheter
och förvaltning av
nätverken,
kommunikation och
publikationer, effekter
på turismen och
ekonomin, finansiell
situation och styrning
Reaktiv övervakning av
hotade platser
Nej
Ja
Nej
Återkallande möjligt
Ja
Ja
Ja, efter ett år av
särskild övervakning
Källa: Revisionsrätten, på grundval av 1) beslut nr 1194/2011/EU om inrättande av Europeiska unionens
insats för det europeiska kulturarvsmärket (EUT L 303, 22.11.2011, s. 1), 2) 2017 års operativa riktlinjer för
genomförandet av Världsarvskonventionen och 3) information från Europarådets kulturvägar och resolution
CM/Res(2013)67 om ändring av reglerna för tilldelning av utmärkelsen ”europeisk kulturväg”.
Bilaga VIII – Utveckling av Eruf-ramen för investeringar i kulturplatser
2007–20131)
2014–20202)
Kommissionens förslag för 2021–2027 3)
Prioriteringar för
investeringar
avseende
kulturplatser
Inga särskilda mål eller
investeringsprioriteringar
fastställdes i
förordningen
Särskilt mål 5 i: ”främja en integrerad social,
ekonomisk och miljömässig utveckling,
kulturarvet och säkerhet i stadsområden”
Särskilt mål 5 ii: ”främja en integrerad, social,
ekonomisk och miljömässig lokal utveckling,
kulturarvet och säkerhet, inklusive på
landsbygden och i kustområden, även genom
lokalt ledd utveckling”
Utgiftskoder
Skydd och bevarande
av kulturarvet
Utveckling av
infrastruktur för kultur,
exklusive kulturella
tjänster
Investeringsprioritering 6c: ”bevara, skydda,
främja och utveckla natur- och kulturarvet”
Investeringsprioritering 8b: ” ökad tillgång till
och utveckling av specifika natur- och
kulturresurser”
Investeringsprioritering 9a: ”investera i
infrastruktur på  det sociala området
genom förbättrad tillgång till sociala och
kulturella tjänster samt rekreationstjänster ”
Outputindikatorer
Ingen kärnindikator
fastställd för
kulturplatser
Resultatindikatorer
Ingen kärnindikator
fastställd för kultur
Skydd, utveckling och främjande av
offentliga kulturtillgångar och kulturarv
Hållbar turism
Ökning av antalet förväntade besök på kulturoch naturarvsplatser och turistattraktioner som
får stöd”
Inga gemensamma resultatindikatorer
fastställdes i förordningen
Skydd, utveckling och främjande av
kulturarv och kulturella tjänster
Gemensam indikator:
RCO 77 – Kapacitet hos kultur- och
turistinfrastruktur som får stöd
Gemensamma indikatorer:
RCR 77 – Antalet turister/besök till platser
som får stöd
RCR 78 – Användare som har nytta av
kulturinfrastruktur som får stöd
Källor: Revisionsrätten, på grundval av följande: 1)Förordning 1083/2006 och förordning 1828/2006. 2)Förordning 1301/2013. 3)Vad beträffar utgiftskoder, se förslaget
till förordning om gemensamma bestämmelser, COM(2018) 375 final, bilagorna 1–22, 29.5.2018; vad beträffar återstående information, se förslaget till förordning
om Europeiska regionala utvecklingsfonden och Sammanhållningsfonden, bilagorna 1 och 2, COM(2018) 372 final, 29.5.2018.
Bilaga IX – Viktigaste målen för insatsområdena i urvalet och mätning av dem med
resultatindikatorer
Sociala
2014–2020
Kulturella
2007–2013
2014–2020
Ekonomiska
2007–2013
2014–2020
2007–2013
Kroatien
Öka sysselsättningen
Resultatindikator
finns trots att mål
inte har fastställts
Förbättra
kulturarvet
Inget mål och ingen
resultatindikator
fastställd
Öka
sysselsättningen
och intäkterna från
turism
Frankrike
Främja social
omvandling
Främja den sociala
sammanhållningen
Bevara och utveckla
det regionala
kulturarvet
Upprusta
kulturarvsplatser och
bygga Louvre-Lensmuseet
Främja ekonomisk
omvandling
Stärka den regionala
spetskompetensen och
attraktionskraften
Tyskland
Inget mål och
ingen resultatindikator har
fastställts
Resultatindikator
finns trots att mål
inte har fastställts
Göra användningen
av kulturarvet
hållbarare
Inget mål och ingen
resultatindikator
fastställd
Bevara städernas
attraktivitet
Utnyttja turismpotentialen
för att öka konkurrenskraften
Italien
Förbättra
villkoren och
reglerna för
användning av
kulturarvet
Förbättra
användningen av
kultur- och
naturresurser
Förbättra villkoren
och reglerna för
utbudet av
kulturarvet
Förbättra bevarandet
av kultur- och
naturresurser
Främja kulturarvet
och turismen för
nationell tillväxt
Öka regionala territoriers
attraktivitet
Utveckla företagsklimatet
och små och medelstora
företags konkurrenskraft
Sociala
Kulturella
Ekonomiska
Polen
Förbättra
tillgängligheten
till
kulturplatser
Öka tillgången till
kultur och använda
kulturarvet
ändamålsenligt
Inget mål och ingen
resultatindikator
fastställd
Förbättra den
kulturella
infrastrukturen och
bevara kulturarvet
Förbättra den
ekonomiska
konkurrenskraften
Öka Polens attraktivitet
Portugal
Öka tillfredsställelsen bland
de boende
Lokal och urban
sammanhållning
genom stärkande av
kollektiva tjänster
Främja stärkande av
kulturarvet
Främja kultur och
kreativitet
Befästa regionen
som en
turistdestination
Ekonomiskt främjande av
specifika resurser
Rumänien
Öka
livskvaliteten
Skapa jobb genom
att utveckla
turismen
Bevara och ta
tillvara kulturarv och
identitet
Restaurering och
hållbart
tillvaratagande av
kulturarv
Stärka den lokala
utvecklingen
Hållbar utveckling och
hållbart främjande av turism
Källa: Revisionsrätten.
Ingen resultatindikator för det målet
Mellan en och två resultatindikatorer
Tre eller fler resultatindikatorer
Akronymer och förkortningar
Eruf: Europeiska regionala utvecklingsfonden.
ESI-fonder: europeiska struktur- och investeringsfonder.
GD: generaldirektorat.
OP: operativt program.
Ordlista
ekonomiskt mål: ett mål som i regel avser produktivitet och/eller sysselsättning.
europeiska struktur- och investeringsfonder (ESI-fonder): de fem viktigaste EUfonderna som tillsammans stöder den ekonomiska utvecklingen i EU, nämligen
Europeiska regionala utvecklingsfonden, Europeiska socialfonden,
Sammanhållningsfonden, Europeiska jordbruksfonden för landsbygdsutveckling och
Europeiska havs- och fiskerifonden; de regleras av en gemensam uppsättning regler.
kulturellt mål: ett mål för att skydda och främja den materiella och immateriella
kulturella mångfalden (kulturplatser, musikframträdanden, konstutställningar etc.).
operativt program: den grundläggande ramen för genomförande av EU-finansierade
sammanhållningsprojekt under en fastställd period som återspeglar de prioriteringar
och mål som fastställts i partnerskapsöverenskommelser mellan kommissionen och
enskilda medlemsstater.
partnerskapsöverenskommelse: en överenskommelse mellan kommissionen och en
medlemsstat eller ett tredjeland/tredjeländer inom ramen för ett av EU:s
utgiftsprogram, i vilken exempelvis strategiska planer, investeringsprioriteringar eller
handelsvillkor eller villkor för tillhandahållande av utvecklingsbistånd fastställs.
socialt mål: ett mål som syftar till att ge alla samhällsgrupper (även missgynnade
personer och personer med funktionsnedsättningar) tillgång till kulturplatser,
demokratisera kunskap och främja utbildning och sysselsättning.
KOMMISSIONENS SVAR PÅ EUROPEISKA REVISIONSRÄTTENS SÄRSKILDA
RAPPORT
EU:S INVESTERINGAR I KULTURPLATSER: ÖKAT FOKUS OCH BÄTTRE
SAMORDNING BEHÖVS”
SAMMANFATTNING
VI: Andra strecksatsen – Den strategiska ramen för kulturpolitiken i Europeiska unionen, utformad av
Europeiska kommissionen (se särskilt En ny europeisk agenda för kultur), är inriktad på kulturens
bidrag till Europas samhällen, ekonomier och internationella förbindelser. Den inriktas inte särskilt på
främjandet av kulturplatser.
Erufs investeringar i restaurering av kulturplatser gör det ofta möjligt för dessa platser att sedan delta i
EU:s kulturinitiativ.
Tredje strecksatsen: Erufs främsta mål är att bidra till att stärka den ekonomiska, sociala och
territoriella sammanhållningen. Enligt punkt 11 i ingressen till Eruf-förordningen bör Eruffinansiering av kultur och stöd till kulturarv grundas på om verksamheten ingår i en territoriell strategi
för ett särskilt område eller i vilken utsträckning den bidrar till sysselsättningsfrämjande tillväxt.
Dessutom är kultur ett område på vilket främst medlemsstaten är behörig, och där Europeiska
kommissionen måste följa subsidiaritetsprincipen.
VII: De ekonomiska och sociala målen för Erufs operativa program och projekt ligger vanligen i linje
med den rättsliga grunden för sammanhållningspolitiken i fördraget.
VIII. a) Kommissionen godtar rekommendationen.
Kommissionen godtar rekommendationen.
Kommissionen godtar rekommendationen.
Redan i omnibusförordningen som trädde i kraft 2018 infördes ytterligare möjligheter till förenklade
kostnadsalternativ för Erufs medfinansiering, och dessa möjligheter utvidgades även i kommissionens
förslag som ska gälla efter 2020.
Enligt kommissionens förslag måste de förvaltande myndigheterna kontrollera att stödmottagarna har
de nödvändiga ekonomiska resurserna och mekanismerna för att täcka drifts- och
underhållskostnader.
Kommissionen godtar rekommendationen.
IAKTTAGELSER
Den strategiska ramen för EU:s åtgärder återspeglar fördragen och EU:s stödjande roll i förhållande
till kultur. Dessutom analyseras i den föreliggande rapporten endast de tillgängliga medlen för
kulturella infrastrukturprojekt (dvs. ESI-fonder), samtidigt som antagandet som görs här rör EUfinansiering totalt sett.
När det gäller Erufs investeringar är målet social och ekonomisk utveckling. Alla investeringar
med en kulturell dimension måste bidra till att uppnå detta mål. Ramen för Erufs stöd anges i bilaga I
till förordningen om gemensamma bestämmelser.
Kommissionen skiljer mellan en EU-ram för investeringar i kulturplatser och en EU-ram för EU:s
åtgärder för kultur.
Det finns bara en strategisk EU-ram för kultur, dvs. den nya europeiska agendan för kultur.
Den enda EU-fond som är särskilt inriktad på kultur är programmet Kreativa Europa, som tar
hänsyn till EU:s aktuella agenda för kultur.
Andra EU-fonder har andra mål och är beroende av andra politiska strategier.
Ingen av de befintliga EU-utmärkelserna för kultur utformades med tanke på att de senare skulle
utlösa EU-finansiering. Kommissionens kulturinitiativ och Eruf-finansiering har skilda mål, och de är
inte avhängiga varandra.
Europeiska kulturarvsmärket och andra kommissionsinitiativ, t.ex. Europeisk kulturhuvudstad,
tilldelas ofta städer/platser som tidigare gynnades av Erufs investeringar. Stödet från Eruf gjorde det
möjligt för dem att därefter få utmärkelsen. Ett bra exempel på detta är Wroclaw, som tack vare Erufs
investeringar under perioden 2007–2013 blev Europeisk kulturhuvudstad 2016.
Fastställandet av kriterier för att välja ut projekt och urvalet ansvarar medlemsstaterna för.
Övervakningskommittén ska granska och godkänna den metod och de kriterier som används för att
välja ut insatser (artikel 110.2a i förordningen om gemensamma bestämmelser).
De olika EU-fonderna är utformade för att komplettera varandra. När det gäller ESI-fonder med
delad förvaltning ska medlemsstaterna fastställa ”Bestämmelser enligt medlemsstaternas
institutionella ramar för samordningen mellan de europeiska struktur- och investeringsfonderna och
andra finansieringsinstrument på unionsnivå och nationell nivå samt med EIB” i partnerskapsavtalen
(artikel 15.1b i i förordningen om gemensamma bestämmelser).
Kravet att inrätta arrangemang som säkerställer samordning mellan ESI-fonderna och andra
finansieringsinstrument på unionsnivå och nationell nivå samt med EIB innebär inte att detaljerade
samordningsmekanismer för varje specifik typ av investeringar som finansieras genom ESI-fonderna
ska upprättas. Detta gäller särskilt investeringar som t.ex. stöd till kulturplatser, som är av begränsad
storlek i de flesta av Erufs program.
Se kommissionens svar på punkt 23.
Enligt förordningen om gemensamma bestämmelser ska medlemsstaterna rapportera ekonomiska
uppgifter till kommissionen på ett systematiskt sätt för Eruf (malltabeller för regelbunden rapportering
anges i kommissionens genomförandeförordning).
Det finns ingen särskild EU-förordning om kulturstatistik. Huvuddelen av EU:s statistik över
kultur härrör från olika undersökningar och datainsamlingar som är reglerade (obligatoriska), t.ex. den
europeiska arbetskraftsundersökningen, statistik över företagsstrukturer och nationalräkenskaper.
Kulturobjekt kan dock inte alltid särskiljas i resultaten från dessa undersökningar (dvs. detaljer som är
relevanta för kultur finns inte tillgängliga i uppgifter som skickas till Eurostat).
Kommissionen erinrar om att Eruf inte är avsett att tillhandahålla sådana ramar för kulturplatser.
Kommissionen betonar att EU inte har behörighet att fastställa ramar för investeringar i kulturplatser,
utan att det är en fråga för medlemsstaterna.
Kommissionen noterar att begränsningen till småskalig kulturell infrastruktur inte var en del av
kommissionens förslag till den nuvarande Eruf-förordningen (COM(2011) 614 final) utan infördes av
medlagstiftarna i förhandlingarna med Europaparlamentet och rådet.
Kommissionen måste prioritera investeringar i kultur jämfört med andra sektorer som transport
eller miljö och se till att förutsättningarna finns för att maximera deras effekter, vilket är orsaken till
att det kan bli vissa minskningar.
Kommissionen betonar att den endast kan kräva att medlemsstaterna utformar sina
partnerskapsöverenskommelser och operativa program i enlighet med de förordningar som godkänts
av medlagstiftarna. Enligt förordningen om gemensamma bestämmelser ska medlemsstaterna använda
ESI-fonder för att på ett effektivt sätt bidra till unionens strategi för smart och hållbar tillväxt för alla.
Det kräver ingen anpassning till någon kulturagenda.
Kommissionen anser att Eruf-investeringarnas ändamålsenlighet endast kan bedömas i förhållande
till Erufs mål, dvs. att främja ekonomisk, social och territoriell sammanhållning.
Fokus för Eruf-finansierade projekt beror på det tematiska mål enligt vilket de finansieras. De
tematiska målen 1–3 inriktas förvisso på tillväxt och konkurrenskraft. Kulturprojekt enligt tematiskt
mål 6 syftade emellertid till att bevara och skydda miljön och främja ett effektivt resursutnyttjande.
Om en investering ägde rum enligt tematiskt mål 9 (t.ex. för tillgång till kulturtjänster) inriktades den
på att främja social delaktighet samt på att bekämpa fattigdom och all diskriminering.
Gemensamt svar 63 och 64
Kommissionen understryker att även om vissa resultatindikatorer inte uppnåddes vid den tidpunkt då
de underliggande projekten avslutades, kan de nås vid tidpunkten då respektive program avslutades,
eftersom det tar tid för resultaten att realiseras.
Kommissionen noterar att det finns lagstiftningskrav för att ange resultatindikatorer för prioriterade
områden, men inte på projektnivå.
Kommissionen betonar att strängare krav för rapportering av resultat har införts i och med
programplaneringsperioden 2014–2020. Revisioner på nationell nivå och på EU-nivå genomförs för
system som används för att samla in, kontrollera och rapportera indikatorer. Otillförlitliga resultat
betraktas som en svaghet i förvaltnings- och kontrollsystemet och kan leda till inställning av
betalningar.
Kommissionen anser att det visserligen fortfarande finns utrymme för förbättringar men att det är
viktiga steg och ett starkt incitament för programmyndigheterna att uppnå ökad tillförlitlighet.
Kommissionen noterar att en delrestaurering i vissa fall var en nödvändighet i den meningen att
underlåtenhet att ingripa kunde ha lett till en stängning av platsen, och därför är det inte alltid ett mål i
sig att öka antalet besökare.
När det gäller Eruf och den gemensamma indikatorn ”ökning av antalet förväntade besök på kulturoch naturarvsplatser” uttrycker denna den förväntade ökningen av antalet besök på en plats året efter
projektets slutförande. De förvaltande myndigheterna fastställer metoden för att uppskatta det
förväntade antalet som kan baseras på efterfrågeanalys. De förvaltande myndigheterna behöver inte
rapportera det faktiska antalet besökare enligt denna gemensamma indikator.
Vid delad förvaltning övervakar kommissionen aggregerade resultat och resultat på program- och
prioriteringsnivå. Det finns inget lagstiftningskrav på att ange resultatindikatorer på projektnivå. En
väl utformad interventionslogik ska säkerställa att utfall och resultat på projektnivå bidrar till att nå de
förväntade resultaten för de operativa programmen, som även de påverkas av externa faktorer. Därför
anser kommissionen att bedömningen av projektens bidrag till programmets mål uttryckt med deras
resultatindikatorer inte kan mätas genom resultatet av enskilda projekt, utan kräver en
konsekvensutvärdering.
Kommissionen delar denna oro och påminner om att det finns en rättslig skyldighet för
stödmottagaren att återbetala EU-bidraget i händelse av en väsentlig förändring av insatsen inom fem
år efter slutbetalningen till stödmottagaren (artikel 71 i förordningen om gemensamma bestämmelser).
I detta avseende kan underlåtenheten att underhålla en restaurerad kulturplats utgöra en väsentlig
förändring av villkoren för insatsens genomförande som underminerar de ursprungliga målen för
Erufs investering.
Tilldelningen av Eruf-medel till projekt drivs av sammanhållningspolitikens mål och av de
särskilda mål som formuleras för de operativa programmen, som oftast inte är kulturinriktade.
Kommissionen betonar att den inte har befogenheter att sträcka sig längre än rapporteringskraven i
artikel 6 i beslut nr 1313/2013/EU om en civilskyddsmekanism för unionen. Detta kräver att
medlemsstaterna ger kommissionen tillgång till en sammanfattning av sina riskbedömningar och en
bedömning av sin riskhanteringsförmåga, med fokus på viktiga risker som fastställts på nationell
(eller regional) nivå.
Den gemensamma indikatorn ”ökningen av antalet besökare på platserna” används endast av de
operativa programmen när det är relevant för de insatser som stöds. Erufs stöd förhindrar inte
nationella myndigheter att vidta åtgärder för bevarande av kulturarv.
Se kommissionens svar på punkt 17.
Denna fråga nämns också i reglerna om undantag från statligt stöd, som måste respekteras från
och med 2014 när Eruf-stöd beviljas. Dessa regler anger särskilt att stödbeloppet för investeringar i
kultur och kulturarv inte får överstiga skillnaden mellan de stödberättigande kostnaderna och
rörelseresultatet för investeringen.
Att resultatindikatorerna för projekt inom Eruf-programmen 2007–2013 inte uppnåddes medförde
inga ekonomiska konsekvenser, eftersom en sådan bestämmelse inte ingick i förordningarna för
2007–2013. Vid delad förvaltning kan de incitamentsmekanismer som Europeiska revisionsrätten
hänvisar till endast tillämpas i avtalsarrangemangen mellan projektstödmottagaren och den
förvaltande myndigheten.
Enligt förordningen om gemensamma bestämmelser ska insatser som medfinansierats av Eruf
upprätthålla sin karaktär, sina mål och genomförandevillkoren under en period på minst fem år från
slutbetalningen till stödmottagaren. Medlemsstaterna övervakar efterlevnaden av denna
lagbestämmelse.
Det nuvarande kravet på utvärdering av effekterna av alla Eruf-insatser utgör ett incitament för
medlemsstaterna att anta ett medellångt perspektiv när de planerar och programplanerar
genomförandet av insatserna, vilket även implicit sörjer för investeringsresultatens varaktighet. Den
direkta övervakningen av varaktigheten hos projektresultaten är dock fortfarande medlemsstaternas
ansvar.
SLUTSATSER OCH REKOMMENDATIONER
Kommissionen noterar att EU:s utmärkelser/initiativ ofta tilldelas de platser som nyligen byggts
eller renoverats tack vare Eruf-finansiering.
Rekommendation 1 – Utforma en lämplig ram för kultur i enlighet med de befogenheter som
anges i fördragen
Kommissionen godtar rekommendationen.
Rekommendation 2 – Se till att privata medel kanaliseras till skyddet av Europas kulturarv
Kommissionen godtar rekommendationen.
Eruf-förordningen behandlar inte fysisk bevarande av finansierade kulturplatser som ett
självständigt mål. Utan att vara en del av en nationell eller regional utvecklingsstrategi kan Eruf
dessutom inte finansiera bevarandet av hotade platser.
Kommissionen noterar att förordningen om gemensamma bestämmelser inte kräver en
övervakning av projektens prestation efter den lagfästa femåriga varaktighetsperioden. Det nuvarande
kravet på utvärdering av effekterna av alla Eruf-insatser utgör ett incitament för medlemsstaterna att
anta ett medellångt perspektiv när de planerar och programplanerar genomförandet av insatserna,
vilket även implicit sörjer för investeringsresultatens varaktighet. Den direkta övervakningen av
varaktigheten hos projektresultaten är dock fortfarande medlemsstaternas ansvar.
Tillämpning av incitaments- och sanktionssystem beroende på projektens prestation faller under
nationell behörighet.
Rekommendation 3 – Stärk den finansiella hållbarheten för kulturplatser som finansieras av
Eruf
Kommissionen godtar rekommendationen.
Redan i omnibusförordningen som trädde i kraft 2018 infördes ytterligare möjligheter till förenklade
kostnadsalternativ för Erufs medfinansiering, och dessa möjligheter utvidgades även i kommissionens
förslag som ska gälla efter 2020.
Enligt kommissionens förslag måste de förvaltande myndigheterna kontrollera att stödmottagarna har
de nödvändiga ekonomiska resurserna och mekanismerna för att täcka drifts- och
underhållskostnader.
Rekommendation 4 – Vidta mer specifika åtgärder för att bevara kulturarvsplatser
Kommissionen godtar rekommendationen.
Granskningsteam
I våra särskilda rapporter redovisar vi resultatet av våra revisioner av EU:s politik och
program eller av förvaltningsteman kopplade till specifika budgetområden. För att
uppnå så stor effekt som möjligt väljer vi ut och utformar granskningsuppgifterna med
hänsyn till riskerna när det gäller prestation eller regelefterlevnad, storleken på de
aktuella intäkterna eller kostnaderna, framtida utveckling och politiskt intresse och
allmänintresse.
Denna effektivitetsrevision utfördes av revisionsrättens avdelning II investeringar för
sammanhållning, tillväxt och inkludering, där ledamoten Iliana Ivanova är ordförande.
Revisionen leddes av revisionsrättens ledamot Pietro Russo med stöd av
Chiara Cipriani (kanslichef), Benjamin Jakob (attaché), Emmanuel Rauch (förstechef),
Sara Pimentel (uppgiftsansvarig) och Ana Popescu, Bernard Witkos,
Dana Smid Foltynova, Jussi Bright, Paulo Manuel Carichas, Sabine Maur-Helmes,
Thierry Lavigne och Tristan Le Guen (revisorer). Hannah Critoph och Richard Moore gav
språkligt stöd.
Från vänster: Sabine Maur-Helmes, Tristan Le Guen, Chiara Cipriani, Benjamin Jakob,
Pietro Russo, Emmanuel Rauch, Sara Pimentel, Jussi Bright och Dana Smid Foltynova.
Tidslinje
Händelse
Revisionsplanen antogs/Revisionen inleddes
Datum
2018
Den preliminära rapporten skickades officiellt till kommissionen
(eller andra revisionsobjekt)
2020
Den slutliga rapporten antogs efter det kontradiktoriska
förfarandet
2020
Kommissionens (eller andra revisionsobjekts) officiella svar
hade tagits emot på alla språk
2020
UPPHOVSRÄTT
© Europeiska unionen 2020.
Europeiska revisionsrättens policy för vidareutnyttjande regleras av Europeiska revisionsrättens beslut
nr 6-2019 om öppen datapolitik och vidareutnyttjande av handlingar.
Om inget annat anges (t.ex. i enskilda meddelanden om upphovsrätt) omfattas revisionsrättens innehåll
som ägs av EU av den internationella licensen Creative Commons Erkännande 4.0 (CC BY 4.0). Det
innebär att vidareutnyttjande är tillåtet under förutsättning att ursprunget anges korrekt och att det
framgår om ändringar har gjorts. Vidareutnyttjas materialet får handlingarnas ursprungliga betydelse
eller budskap inte förvanskas. Revisionsrätten bär inte ansvaret för eventuella konsekvenser av
vidareutnyttjande.
När enskilda privatpersoner kan identifieras i ett specifikt sammanhang, exempelvis på bilder av
revisionsrättens personal, eller om arbete av tredje part används, måste tillstånd inhämtas med
avseende på de ytterligare rättigheterna. Om tillstånd beviljas upphävs det allmänna godkännande som
nämns ovan, och eventuella begränsningar av materialets användning måste tydligt anges.
För användning eller återgivning av innehåll som inte ägs av EU kan tillstånd behöva inhämtas direkt från
upphovsrättsinnehavarna.
Foto ruta 1: © Capital Europeia da Cultura Guimarães 2012.
Bild 2: Ikoner gjorda av Pixel perfect från https://flaticon.com.
Foton ruta 3: © Katowices stad.
Foto ruta 4: © Fotograf: Luciano Romano.
Foto ruta 7: © Fotograf: Henrique Patricio.
Foto 1 ruta 10: Källa: Scheda ispettiva, Casa dell’Efebo I 7, 11, från Parco Archeologico di Pompei.
Foto 2 ruta 10: Källa: Relazione tecnica, Casa dell’Efebo, januari 2016, från Parco Archeologico di
Pompei.
Programvara eller handlingar som omfattas av immateriella rättigheter, till exempel patent,
varumärkesskydd, mönsterskydd samt upphovsrätt till logotyper eller namn, omfattas inte av
revisionsrättens policy för vidareutnyttjande eller av licensen.
EU-institutionernas webbplatser inom domänen europa.eu innehåller länkar till webbplatser utanför
den domänen. Eftersom revisionsrätten inte kontrollerar dem uppmanas du att ta reda på vilken
integritets- och upphovsrättspolicy de tillämpar.
Användning av Europeiska revisionsrättens logotyp
Europeiska revisionsrättens logotyp får inte användas utan Europeiska revisionsrättens
förhandsgodkännande.
PDF
HTML
ISBN 978-92-847-4442-8 ISSN 1977-5830
ISBN 978-92-847-4461-9 ISSN 1977-5830
doi:10.2865/8369
doi:10.2865/584843
QJ-AB-20-005-SV-N
QJ-AB-20-005-SV-Q
På kulturområdet fastställer fördraget som överordnat mål att EU
ska respektera rikedomen hos sin kulturella mångfald och sörja
för att det europeiska kulturarvet skyddas och utvecklas.
Eftersom kulturfrågor huvudsakligen är medlemsstaternas
behörighet kan unionen endast uppmuntra till samarbete mellan
medlemsstater och stödja eller komplettera deras insatser.
Vi bedömde de ekonomiska, sociala och kulturella effekterna av
Eruf-investeringar i kulturplatser och kulturplatsernas finansiella
och fysiska hållbarhet. Vi granskade kommissionens arbete och
bedömde 27 projekt i sju medlemsstater.
Slutsatsen av revisionen är att den nuvarande ramen saknar fokus
och behöver samordnas bättre för att säkerställa att Erufinvesteringarna i kulturplatser blir ändamålsenliga och hållbara.
Revisionsrättens särskilda rapport i enlighet med artikel 287.4
andra stycket i EUF-fördraget.
