SKLEP SODIŠČA (tretji senat)
z dne 17. januarja 2012(*)
Avtorska pravica – Informacijska družba – Direktiva 2001/29/ES – Člen 5(1) in (5) – Književna in umetniška dela – Reproduciranje kratkih odlomkov književnih del – Časopisni članki – Začasno in prehodno reproduciranje – Tehnološki proces, ki zajema skeniranje člankov s poznejšo pretvorbo v tekstovno datoteko, elektronsko obdelavo reprodukcije ter shranjevanje dela te reprodukcije – Začasna dejanja reproduciranja, ki so sestavni in bistveni del takega tehnološkega procesa – Namen teh dejanj, ki je zakonita uporaba zaščitenega dela ali predmeta sorodnih pravic – Neodvisni ekonomski pomen navedenih dejanj“
V zadevi C‑302/10,
katere predmet je predlog za sprejetje predhodne odločbe na podlagi člena 267 PDEU, ki ga je vložilo Højesteret (Danska) z odločbo z dne 16. junija 2010, ki je prispela na Sodišče 18. junija 2010, v postopku
Infopaq International A/S
proti
Danske Dagblades Forening,
SODIŠČE (tretji senat),
v sestavi K. Lenaerts, predsednik senata, J. Malenovský (poročevalec), E. Juhász, G. Arestis in T. von Danwitz, sodniki,
generalna pravobranilka: V. Trstenjak,
sodni tajnik: A. Calot Escobar,
na podlagi pisnega postopka,
ob upoštevanju stališč, ki so jih predložili:
za Infopaq International A/S A. Jensen, odvetnik,
za Danske Dagblades Forening M. Dahl Pedersen, odvetnik,
za špansko vlado N. Díaz Abad, zastopnica,
za Evropsko komisijo J. Samnadda in H. Støvlbæk, zastopnika,
po odločitvi Sodišča, da odloči z obrazloženim sklepom v skladu s členom 104(3), prvi pododstavek, Poslovnika,
sprejema naslednji
Sklep
Predlog za sprejetje predhodne odločbe se nanaša na razlago člena 5(1) in (5) Direktive 2001/29/ES Evropskega parlamenta in Sveta z dne 22. maja 2001 o usklajevanju določenih vidikov avtorske in sorodnih pravic v informacijski družbi (UL, posebna izdaja v slovenščini, poglavje 17, zvezek 1, str. 230).
Ta predlog je bil vložen v okviru spora med družbo Infopaq International A/S (v nadaljevanju: Infopaq) in združenjem Danske Dagblades Forening (v nadaljevanju: DDF) glede zavrnitve zahtevka družbe Infopaq za priznanje, da ji ni bilo treba pridobiti privolitve imetnikov avtorskih pravic za dejanja reproduciranja časopisnih člankov z avtomatiziranim procesom, ki zajema njihovo skeniranje in pretvorbo v digitalno datoteko s poznejšo elektronsko obdelavo te datoteke.
Pravni okvir
Pravo Unije
V uvodnih izjavah 4, od 9 do 11, 21, 22, 31 in 33 Direktive 2001/29 je navedeno:
Usklajena pravna ureditev avtorske in sorodnih pravic bo zaradi večje pravne varnosti in hkrati z zagotavljanjem visoke stopnje varstva intelektualne lastnine omogočala naložbe v ustvarjalnost in inovacije vključno z omrežno infrastrukturo
Vsakršno usklajevanje avtorske in sorodnih pravic mora temeljiti na visoki stopnji varstva, kajti takšne pravice so za intelektualno ustvarjanje bistvenega pomena.
Če naj avtorji ali izvajalci nadaljujejo z ustvarjalnim in umetniškim delom, morajo za uporabo svojega dela prejeti primerno nagrado
Dodano je, da je strog, učinkovit sistem varstva avtorske in sorodnih pravic eden glavnih načinov za zagotavljanje, da evropska kulturna ustvarjalnost in proizvodnja prejmeta nujna sredstva ter za varovanje neodvisnosti in dostojanstva umetniških ustvarjalcev in izvajalcev.
Ta direktiva naj določi obseg dejanj, ki jih zajema pravica reproduciranja za različne upravičence. To naj poteka v skladu s pravnim redom Skupnosti. Potrebna je široka opredelitev teh dejanj, ki bo zagotovila pravno varnost na notranjem trgu.
Cilja ustrezne podpore razširjanju kulture se ne sme doseči z žrtvovanjem strogega varstva pravic ali z dopuščanjem nezakonitih oblik distribuiranja ponarejenih ali piratskih del.
Zagotoviti je treba pravično ravnotežje pravic in interesov med različnimi kategorijami imetnikov pravic, pa tudi med različnimi kategorijami imetnikov pravic in uporabnikov varovanih predmetov.
Izključna pravica reproduciranja naj ima izjemo, ki naj dopušča določena dejanja začasnega reproduciranja, ki so prehodne ali naključne reprodukcije in so sestavni in nujni del tehnološkega procesa ter se izvajajo zgolj zato, da se omogoči bodisi učinkovit prenos v omrežju med tretjimi strankami preko posrednika bodisi zakonita uporaba dela ali predmeta. Takšna dejanja reproduciranja ne smejo imeti lastne ekonomske vrednosti. Kolikor ustrezajo tem pogojem, naj ta izjema zajema dejanja, ki omogočajo brskanje, pa tudi dejanja predpomnjenja vključno s tistimi, ki omogočajo učinkovito delovanje prenosnih sistemov, pod pogojem, da vmesnik ne spreminja informacij in se ne vmešava v zakonito uporabo tehnologije, ki jo široko priznava in uporablja industrija, za pridobivanje podatkov o uporabi informacij. Uporaba velja za pravilno, kadar je odobrena s strani imetnika pravic oziroma kadar je ne omejuje zakon.“
Člen 1(1) Direktive 2001/29 določa:
Ta direktiva ureja pravno varstvo avtorske in sorodnih pravic v okviru notranjega trga s posebnim poudarkom na informacijski družbi.“
Člen 2(a) te direktive določa:
Države članice predvidijo za spodaj naštete izključno pravico, da dovolijo ali prepovedo, neposredno ali posredno, začasno ali stalno, reproduciranje na vsak način in v vsaki obliki, v celoti ali deloma:
avtorjem za njihova dela“.
Člen 5 navedene direktive določa:
Začasna dejanja razmnoževanja [reproduciranja] iz člena 2, ki so prehodna ali spremljevalna ter so sestavni in bistveni del tehnološkega procesa in katerih edini namen je omogočiti:
prenos po omrežju med tretjimi strankami po posredniku, ali
zakonito uporabo
dela ali predmeta sorodnih pravic, ki naj se izvede in ki nima nobenega neodvisnega ekonomskega pomena, so izvzeta iz pravice reproduciranja, ki jo določa člen 2.
Države članice lahko predvidijo izjeme in omejitve pravic iz členov 2 in 3 v naslednjih primerih:
reproduciranje v tisku, priobčitev javnosti oziroma dajanje na voljo javnosti objavljenih člankov o aktualnih gospodarskih, političnih ali verskih temah oziroma predvajanih del ali druge vsebine istega značaja v primerih, ko takšna uporaba ni izrecno prepovedana in dokler je naveden vir vključno z avtorjevim imenom, oziroma uporaba del ali predmetov sorodnih pravic v zvezi s poročanjem o aktualnih dogodkih v obsegu, ki ga upravičuje informativni namen, in ob navedbi vira vključno z avtorjevim imenom, razen če se to izkaže za nemogoče;
citati z namenom kritike ali ocene pod pogojem, da se nanašajo na delo ali na predmet sorodnih pravic, ki je bil že bil zakonito dan na voljo javnosti, da je naveden vir vključno z avtorjevim imenom, razen če se to izkaže za nemogoče, in da je njihova uporaba v skladu s pošteno prakso ter v obsegu, ki ga zahteva poseben namen;
Izjeme in omejitve iz odstavkov 1, 2, 3 in 4 naj se uporabijo le v določenih posebnih primerih, ki niso v nasprotju z normalnim izkoriščanjem dela ali drugega predmeta in ne vplivajo pretirano na legitimne interese imetnika pravic.“
Nacionalno pravo
Člena 2 in 5(1) Direktive 2001/29 sta bila v danski pravni red prenesena s členoma 2 in 11a(1) zakona št. 395 o avtorski pravici (lov n° 395 om ophavsret) z dne 14. junija 1995 (Lovtidende 1995 A, str. 1796), kakor je bil spremenjen in kodificiran med drugim z zakonom št. 1051 (lov n° 1051) z dne 17. decembra 2002 (Lovtidende 2002 A, str. 7881).
Spor o glavni stvari in vprašanja za predhodno odločanje
Družba Infopaq opravlja dejavnosti glede spremljanja in analize tiskanih medijev, ki v bistvu zajemajo pripravljanje povzetkov izbranih člankov iz danskega dnevnega tiska in različnih revij. Ta izbor člankov se opravi glede na teme, ki jih izberejo stranke, v procesu, imenovanem zbiranje podatkov“. Povzetki se pošljejo strankam po elektronski pošti.
Združenje DDF je poklicno združenje danskih dnevnih časopisov, katerega namen je med drugim pomagati članom pri vseh vprašanjih v zvezi z avtorsko pravico.
Združenje DDF je bilo leta 2005 seznanjeno s tem, da družba Infopaq za gospodarske namene obdeluje časopisne članke brez privolitve imetnikov avtorskih pravic na teh člankih. Ker je združenje DDF menilo, da je taka privolitev nujna za obdelavo člankov v zadevnem procesu, je o tem obvestila družbo Infopaq.
Proces zbiranja podatkov ima pet zaporednih faz, ki po mnenju združenja DDF povzročijo štiri dejanja reproduciranja časopisnih člankov.
Prvič, sodelavci družbe Infopaq ročno vpišejo zadevne publikacije v elektronsko bazo podatkov.
Drugič, potem ko se odreže hrbtna stran, se te publikacije skenirajo, tako da so listi med seboj ločeni. Del publikacije, ki bo obdelan, se izbere iz baze podatkov, preden se publikacija vstavi v optični čitalec (skener). Skeniranje omogoča, da se iz vsake strani publikacije ustvari datoteka v obliki TIFF (Tagged Image File Format“, v nadaljevanju: datoteka TIFF). Po koncu tega postopka se datoteka TIFF prenese na strežnik OCR (Optical Character Recognition“) (optično prepoznavanje znakov).
Tretjič, ta strežnik OCR datoteko TIFF pretvori v podatke, ki se lahko računalniško obdelajo. Med tem procesom se slika vsakega znaka spremeni v digitalno kodo, iz katere računalnik razbere vrsto znaka. Na primer, slika črk TDC“ se preoblikuje v podatek, ki ga računalnik lahko obdela kot črke TDC“ in spremeni v tekstovno obliko, ki jo računalniški sistem lahko prepozna. Ti podatki se shranijo kot tekstovne datoteke, ki se lahko preberejo s katerim koli urejevalnikom besedila (v nadaljevanju: tekstovna datoteka). Proces OCR se konča z izbrisom datoteke TIFF.
Četrtič, tekstovna datoteka se analizira, da bi se v njej poiskale predhodno določene ključne besede. Za vsako najdeno besedo se ustvari datoteka, v kateri se navedejo naslov, oddelek in stran publikacije, na kateri je navedena ključna beseda, ter vrednost, izražena v odstotkih od 0 do 100, da bi se označil položaj te ključne besede v besedilu in tako olajšalo branje članka. Da bi se pri branju članka še bolj olajšalo iskanje ključne besede, se skupaj z njo navede še pet besed pred njo in pet besed za njo (v nadaljevanju: odlomek, sestavljen iz enajstih besed). Ta proces se konča z izbrisom tekstovne datoteke.
Petič, proces zbiranja podatkov se konča z izdajo spremnega lista za vsako stran publikacije, na kateri je navedena ključna beseda. Spremni list je lahko na primer tak:
november 2005 – Dagbladet Arbejderen, stran 3:
TDC: 73 % ‚prihodnja prodaja telekomunikacijske skupine TDC, ki bo po pričakovanjih prevzeta‘“.
Družba Infopaq je izpodbijala, da je za tako dejavnost potrebna privolitev imetnikov avtorskih pravic, in je pri Østre Landsret proti združenju DDF vložila tožbo, s katero je predlagala, naj se mu naloži, da družbi Infopaq prizna pravico uporabe zgoraj navedenega procesa brez privolitve tega poklicnega združenja ali njegovih članov. Ker je Østre Landsret to tožbo zavrnilo, je družba Infopaq pri predložitvenem sodišču vložila pritožbo.
Predložitveno sodišče meni, da ni sporno, da privolitev imetnikov avtorskih pravic za opravljanje dejavnosti spremljanja tiskanih medijev in pripravljanja povzetkov ni potrebna, če ta obsega fizično branje vsake publikacije, izbor upoštevnih člankov na podlagi predhodno določenih ključnih besed in ročno izdelavo spremnega lista za avtorja povzetka, na katerem sta navedena ključna beseda v članku in položaj članka v publikaciji. Stranki v postopku v glavni stvari prav tako soglašata glede dejstva, da je pripravljanje povzetka samo po sebi zakonito in da se zanj ne zahteva privolitev imetnikov navedenih pravic.
Poleg tega se ne izpodbija, da navedeni proces zbiranja podatkov vključuje dve dejanji reproduciranja, in sicer izdelavo datotek TIFF pri skeniranju natisnjenih člankov in izdelavo tekstovnih datotek s pretvorbo datotek TIFF. Poleg tega ni sporno, da se pri tem procesu reproducirajo deli skeniranih člankov, saj se odlomek iz enajstih besed shrani v računalniški spomin, enajst besed pa se natisne na papir.
Vendar stranki v postopku v glavni stvari ne soglašata glede vprašanja, ali gre pri zgoraj navedenih dejanjih za dejanji reproduciranja v smislu člena 2 Direktive 2001/29. Prav tako si nasprotujeta glede vprašanja, ali so vsa dejanja v postopku v glavni stvari v tem primeru zajeta z izvzetjem iz pravice reproduciranja, ki ga določa člen 5(1) te direktive.
V teh okoliščinah je Højesteret 21. decembra 2007 prekinilo odločanje in Sodišču v predhodno odločanje predložilo trinajst vprašanj, ki se nanašajo na razlago členov 2(a) ter 5(1) in (5) navedene direktive.
Sodišče je na ta vprašanja odgovorilo s sodbo z dne 16. julija 2009 v zadevi Infopaq International (C‑5/08, ZOdl., str. I‑6569), v kateri je razsodilo, po eni strani, da pojem delnega reproduciranja v smislu člena 2 Direktive 2001/29 lahko zajema dejanje v procesu zbiranja podatkov, in sicer shranjevanje odlomka zaščitenega dela, sestavljenega iz enajstih besed, v računalniški spomin in njegovo tiskanje, če so tako reproducirani elementi lastna intelektualna stvaritev njihovega avtorja, kar mora preveriti predložitveno sodišče. Po drugi strani je Sodišče ugotovilo, da čeprav je člen 5(1) te direktive omogočal izvzetje iz pravice reproduciranja dejanj reproduciranja, ki so prehodna ali spremljevalna, zadnje dejanje v procesu zbiranja podatkov v postopku v glavni stvari, med katerim je družba Infopaq natisnila odlomke, sestavljene iz enajstih besed, ni bilo prehodno ali spremljevalno dejanje. Zato je Sodišče odločilo, da tega dejanja in procesa zbiranja podatkov, katerega del je bilo to dejanje, ni bilo mogoče izvesti brez privolitve imetnikov avtorskih pravic.
Højesteret pa je po tej sodbi ugotovilo, da je lahko še vedno pozvano, naj odloči o tem, ali je družba Infopaq kršila Direktivo 2001/29 z izvedbo navedenega procesa, razen tiska odlomka, sestavljenega iz enajstih besed, in sicer če bi se omejila na izvedbo prvih treh dejanj reproduciranja. Zato se je Højesteret odločilo Sodišču v predhodno odločanje predložiti ta vprašanja:
Ali je stopnja tehnološkega procesa, na kateri se opravi začasno dejanje reproduciranja, pomembna pri ugotavljanju, ali je mogoče to dejanje šteti za ‚sestavni in bistveni del tehnološkega procesa‘ [v smislu člena 5(1) Direktive 2001/29]?
Ali se dejanje reproduciranja lahko šteje za ‚sestavni in bistveni del tehnološkega procesa‘, če zajema ročno skeniranje celotnih časopisnih člankov, s čimer so ti preoblikovani iz tiskanega medija v digitalni medij?
Ali pojem ‚zakonita uporaba‘ iz člena 5(1) Direktive 2001/29 zajema vsako vrsto uporabe, za katero ni potrebna privolitev imetnika avtorskih pravic?
Ali ‚zakonita uporaba‘ iz člena 5(1) Direktive 2001/29 zajema skeniranje celotnih časopisnih člankov, ki ga opravi podjetje, in poznejšo obdelavo reprodukcije za uporabo pri pripravljanju povzetkov, čeprav imetnik avtorskih pravic v ta dejanja ni privolil, če so izpolnjene zahteve iz te določbe?
Ali je za odgovor na to vprašanje pomembno, da se po končanem procesu zbiranja podatkov shrani enajst besed?
Katera merila je treba uporabiti za presojo, ali imajo začasna dejanja reproduciranja ‚neodvisen ekonomski pomen‘ v smislu člena 5(1) Direktive 2001/29, če so izpolnjene druge zahteve iz te določbe?
Ali je mogoče povečanje uporabnikove učinkovitosti zaradi začasnih dejanj reproduciranja upoštevati pri presoji, ali imajo dejanja ‚neodvisen ekonomski pomen‘ v smislu člena 5(1) Direktive 2001/29‘?
Ali se skeniranje celotnih časopisnih člankov, ki ga opravi podjetje, in poznejša obdelava reprodukcije lahko štejeta za ‚določene posebne primere, ki niso v nasprotju z normalnim izkoriščanjem‘ navedenih člankov in ‚ne vplivajo pretirano na legitimne interese imetnika pravic‘ v smislu člena 5(5) Direktive 2001/29, če so izpolnjeni pogoji iz odstavka 1 tega člena?
Ali je za odgovor na to vprašanje pomembno, da se po končanem procesu zbiranja podatkov shrani enajst besed?“
Vprašanja za predhodno odločanje
Sodišče lahko na podlagi člena 104(3), prvi pododstavek, Poslovnika, če je iz obstoječe sodne prakse mogoče jasno sklepati, kakšen bo odgovor na predloženo vprašanje, po opredelitvi generalnega pravobranilca kadar koli odloči z obrazloženim sklepom, v katerem navede ustrezno sodno prakso. To velja v tej zadevi.
Uvodne ugotovitve
Člen 5(1) Direktive 2001/29 določa, da je dejanje reproduciranja izvzeto iz pravice reproduciranja, ki jo določa člen 2 te direktive, le če izpolnjuje pet pogojev, in sicer če je to dejanje:
začasno;
prehodno ali spremljevalno;
sestavni in bistveni del tehnološkega procesa;
če je edini namen tega procesa omogočiti prenos po omrežju med tretjimi strankami po posredniku ali zakonito uporabo dela ali predmeta sorodnih pravic in
če nima nobenega neodvisnega ekonomskega pomena.
Po eni strani je treba spomniti, da so ti pogoji kumulativni, tako da če eden od njih ni izpolnjen, dejanje reproduciranja na podlagi člena 5(1) Direktive 2001/29 ni izvzeto iz pravice reproduciranja, ki jo določa člen 2 te direktive (zgoraj navedena sodba Infopaq International, točka 55).
Po drugi strani je iz sodne prakse Sodišča razvidno, da je treba zgoraj navedene pogoje razlagati ozko, ker člen 5(1) te direktive pomeni izjemo od splošnega pravila, ki ga ta uvaja in ki zahteva, da imetnik avtorske pravice dovoli kakršno koli reproduciranje svojega zaščitenega dela (glej zgoraj navedeno sodbo Infopaq International, točki 56 in 57, in sodbo z dne 4. oktobra 2011 v združenih zadevah Football Association Premier League in drugi, C‑403/08 in C‑429/08, ZOdl., str. I‑9083, točka 162).
V teh okoliščinah je treba preizkusiti vprašanja za predhodno odločanje, s katerimi predložitveno sodišče želi izvedeti, ali dejanja reproduciranja, ki se opravijo med tehničnim procesom, kot je ta v postopku v glavni stvari, izpolnjujejo tretji, četrti in peti pogoj iz člena 5(1) Direktive 2001/29 in pogoje iz člena 5(5) te direktive. Predlog za sprejetje predhodne odločbe pa se ne nanaša na prvi in drugi pogoj iz člena 5(1) navedene direktive, ker je Sodišče o teh pogojih že odločilo v točkah od 61 do 71 zgoraj navedene sodbe Infopaq International.
Prvo in drugo vprašanje v zvezi s pogojem, v skladu s katerim morajo biti dejanja reproduciranja sestavni in bistveni del tehnološkega procesa
Predložitveno sodišče s prvim in drugim vprašanjem, ki ju je treba obravnavati skupaj, v bistvu sprašuje, ali je treba člen 5(1) Direktive 2001/29 razlagati tako, da začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, izpolnjujejo pogoj, v skladu s katerim morajo biti ta dejanja sestavni in bistveni del tehnološkega procesa. V zvezi s tem zlasti sprašuje, ali je treba upoštevati stopnjo tehnološkega procesa, na kateri se ta dejanja opravijo, in to, da navedeni tehnični proces zahteva človeško posredovanje.
Pojem sestavni in bistveni del tehnološkega procesa“ zahteva, da se začasna dejanja reproduciranja opravijo v celoti v okviru izvedbe tehnološkega procesa in da se torej ne opravijo v celoti ali deloma zunaj takega procesa. Ta pojem prav tako predpostavlja, da je izvedba začasnega dejanja reproduciranja nujno potrebna za dobro in učinkovito delovanje tehnološkega procesa (glej v tem smislu zgoraj navedeno sodbo Infopaq International, točka 61).
Poleg tega, ker v členu 5(1) Direktive 2001/29 ni pojasnjeno, na kateri stopnji tehnološkega procesa se morajo opraviti začasna dejanja reproduciranja, ni izključeno, da se s takim dejanjem začne ali konča ta proces.
Prav tako nič v tej določbi ne kaže na to, da tehnološki proces ne sme vključevati nobenega človeškega posredovanja in zlasti da je izključen ročni začetek tega procesa, da bi bila izvedena prva začasna reprodukcija.
V obravnavanem primeru je treba spomniti, da zadevni tehnični proces zajema elektronsko in samodejno iskanje po časopisnih člankih ter ugotavljanje in pridobivanje iz njih predhodno določenih ključnih besed za izboljšanje učinkovitosti priprave povzetkov časopisnih člankov.
V tem okviru se tri dejanja reproduciranja opravijo zaporedoma. Najprej se izdela datoteka TIFF, nato tekstovna datoteka in nazadnje datoteka, ki vsebuje odlomek iz enajstih besed.
Najprej, v zvezi s tem ni sporno, da se nobeno od teh dejanj ne opravi zunaj navedenega tehničnega procesa.
Dalje, ob upoštevanju ugotovitev iz točk od 30 do 32 tega sklepa ni upoštevno, da se tak tehnični proces začne z ročno vstavitvijo časopisnih člankov v optični čitalec s ciljem prve začasne reprodukcije – izdelava datoteke TIFF – in da se konča z začasnim dejanjem reproduciranja, in sicer izdelavo datoteke, ki vsebuje odlomek iz enajstih besed.
Nazadnje je treba poudariti, da so zadevna začasna dejanja reproduciranja nujno potrebna za dobro in učinkovito delovanje zadevnega tehnološkega procesa. Njegov namen je namreč iz časopisnih člankov ugotoviti in izvleči, v digitalni obliki, predhodno določene ključne besede, tako da tako elektronsko iskanje zahteva spremembo teh člankov iz papirne oblike v digitalne podatke, saj je taka sprememba potrebna za prepoznavo navedenih podatkov, za ugotovitev ključnih besed in za to, da se te besede izvleče.
V nasprotju s tem, kar trdi združenje DDF, te ugotovitve ni mogoče izpodbiti s tem, da bi bilo mogoče povzetke časopisnih člankov pripraviti brez reproduciranja. V zvezi s tem zadostuje ugotoviti, da se tak povzetek pripravi zunaj navedenega procesa, saj se opravi za njim in zato ni pomemben za presojo, ali tak proces deluje dobro in učinkovito brez zadevnih dejanj reproduciranja.
Glede na vse navedeno je treba na prvo in drugo vprašanje odgovoriti, da je treba člen 5(1) Direktive 2001/29 razlagati tako, da začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, izpolnjujejo pogoj, v skladu s katerim morajo biti ta dejanja sestavni in bistveni del tehnološkega procesa, ne glede na to, da pomenijo začetek in konec tega procesa ter zahtevajo človeško posredovanje.
Tretje in četrto vprašanje v zvezi s pogojem, v skladu s katerim morajo imeti dejanja reproduciranja samo en namen, in sicer omogočiti bodisi prenos zaščitenega dela ali predmeta sorodnih pravic v omrežju med tretjimi strankami prek posrednika bodisi zakonito uporabo takega dela ali predmeta sorodnih pravic
Predložitveno sodišče s tretjim in četrtim vprašanjem, ki ju je treba obravnavati skupaj, v bistvu sprašuje, ali je treba člen 5(1) Direktive 2001/79 razlagati tako, da so začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, skladna s pogojem, v skladu s katerim morajo imeti dejanja reproduciranja samo en namen, in sicer omogočiti bodisi učinkovit prenos zaščitenega dela ali predmeta sorodnih pravic v omrežju med tretjimi strankami prek posrednika bodisi zakonito uporabo takega dela ali predmeta sorodnih pravic.
Najprej je treba poudariti, da namen zadevnih dejanj reproduciranja ni omogočiti prenos v omrežju med tretjimi strankami prek posrednika. V teh okoliščinah je treba presoditi, ali je edini cilj teh dejanj omogočiti zakonito uporabo zaščitenega dela ali predmeta sorodnih pravic.
V zvezi s tem, kot je razvidno iz uvodne izjave 33 Direktive 2001/29, se uporaba šteje za zakonito, kadar jo je odobril zadevni imetnik pravic ali kadar je ne omejuje veljaven zakon (zgoraj navedena sodba Football Association Premier League in drugi, točka 168).
V zadevi v postopku v glavni stvari je treba po eni strani poudariti, da je v položaju, na katerega se sklicuje predložitveno sodišče, v katerem je bilo zadnje dejanje tehničnega procesa zbiranja podatkov opuščeno, in sicer tisk odlomka, sestavljenega iz enajstih besed, namen zadevnega tehničnega procesa, in zato izdelave datoteke TIFF, tekstovne datoteke in datoteke, ki vsebuje odlomek, sestavljen iz enajstih besed, omogočiti učinkovitejšo pripravo povzetkov časopisnih člankov in s tem njihovo uporabo. Po drugi strani v spisu, predloženemu Sodišču, nič ne kaže na to, da naj bi bil namen rezultata tega tehničnega procesa, in sicer odlomek, sestavljen iz enajstih besed, omogočiti drugačno uporabo.
Glede zakonitosti navedene uporabe ni sporno, da priprave povzetka časopisnih člankov v obravnavani zadevi imetniki avtorskih pravic na teh člankih niso odobrili. Glede na to je treba poudariti, da taka dejavnost ni omejena z zakonodajo Unije. Poleg tega je iz usklajenih izjav družbe Infopaq in združenja DDF razvidno, da priprava navedenega povzetka ni dejavnost, ki je omejena z dansko zakonodajo.
V teh okoliščinah ni mogoče šteti, da je navedena uporaba nezakonita.
Glede na navedeno je treba na tretje in četrto vprašanje odgovoriti, da je treba člen 5(1) Direktive 2001/29 razlagati tako, da so začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, skladna s pogojem, v skladu s katerim morajo imeti dejanja reproduciranja samo en namen, in sicer omogočiti zakonito uporabo dela ali predmeta sorodnih pravic.
Peto in šesto vprašanje v zvezi s pogojem, v skladu s katerim dejanja reproduciranja ne smejo imeti neodvisnega ekonomskega pomena
Ob upoštevanju okvira zadeve v postopku v glavni stvari, kot tudi obsega prejšnjih vprašanj, je treba peto in šesto vprašanje razumeti tako, da se z njima želi izvedeti, ali začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, izpolnjujejo pogoj iz člena 5(1) Direktive 2001/29, v skladu s katerim ta dejanja ne smejo imeti neodvisnega ekonomskega pomena.
V zvezi s tem je treba spomniti, da je namen začasnih dejanj reproduciranja v smislu člena 5(1) omogočiti dostop do zaščitenih del in njihovo uporabo. Ker imajo ta lastno ekonomsko vrednost, imata dostop do njih in njihova uporaba nujno ekonomski pomen (glej v tem smislu zgoraj navedeno sodbo Football Association Premier League in drugi, točka 174).
Poleg tega, kot je razvidno iz uvodne izjave 33 Direktive 2001/29, je namen začasnih dejanj reproduciranja – v tej zadevi dejanj, ki omogočajo brskanje in predpomnenje – olajšati uporabo dela ali izboljšati učinkovitost te uporabe. Tako je s temi dejanji neločljivo povezano povečanje učinkovitosti v okviru take uporabe in zato povečanje dobička ali zmanjšanje stroškov proizvodnje.
Glede na to navedena dejanja ne smejo imeti neodvisnega ekonomskega pomena, kar pomeni, da ekonomske koristi v zvezi z njihovim izvajanjem ne smejo biti niti ločene niti ločljive od ekonomskih koristi v zvezi z zakonito uporabo zadevnega dela, in ne smejo ustvarjati dodatnih ekonomskih koristi, ki presegajo tiste v zvezi z navedeno uporabo zaščitenega dela (glej v tem smislu zgoraj navedeno sodbo Football Association Premier League in drugi, točka 175).
Povečanje učinkovitosti zaradi izvedbe začasnih dejanj reproduciranja, kot so ta v postopku v glavni stvari, nima takega neodvisnega ekonomskega pomena, če se ekonomske koristi v zvezi z njegovo uporabo pojavijo le ob uporabi reproduciranega predmeta, tako da ni niti ločeno niti ločljivo od ekonomskih koristi v zvezi z njegovo uporabo.
V nasprotju s tem so koristi v zvezi z začasnim dejanjem reproduciranja ločene in ločljive, če lahko avtor tega dejanja ustvari dobiček zaradi gospodarskega izkoriščanja samih začasnih reprodukcij.
Enako velja, če začasna dejanja reproduciranja privedejo do spremembe reproduciranega predmeta, kot obstaja ob sprožitvi zadevnega tehničnega procesa, ker namen navedenih aktov ni več olajšati njegovo uporabo, temveč uporabo drugačnega predmeta.
Zato je treba na peto in šesto vprašanje odgovoriti, da je treba člen 5(1) Direktive 2001/29 razlagati tako, da začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, izpolnjujejo pogoj, v skladu s katerim ta dejanja ne smejo imeti neodvisnega ekonomskega pomena, če izvedba teh dejanj ne omogoča ustvarjanja dodatnega dobička, ki presega dobiček v zvezi z zakonito uporabo zaščitenega dela, in če začasna dejanja reproduciranja ne privedejo do spremembe tega dela.
Sedmo vprašanje v zvezi s pogojem, v skladu s katerim dejanja reproduciranja ne smejo biti v nasprotju z običajno uporabo dela in tudi ne smejo nerazumno posegati v zakonite interese imetnika pravic
Predložitveno sodišče s sedmim vprašanjem v bistvu sprašuje, ali je treba člen 5(5) Direktive 2001/29 razlagati tako, da začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, izpolnjujejo pogoj, v skladu s katerim ne smejo biti v nasprotju z običajno uporabo dela in tudi ne smejo nerazumno posegati v zakonite interese imetnika pravic.
V zvezi s tem zadošča ugotoviti, da če ta dejanja reproduciranja izpolnjujejo vse pogoje iz člena 5(1) Direktive 2001/29, kakor so razloženi v sodni praksi Sodišča, je treba šteti, da niso v nasprotju z običajno uporabo dela in tudi nerazumno ne posegajo v zakonite interese imetnika pravic (glej zgoraj navedeno sodbo Football Association Premier League in drugi, točka 181).
Zato je treba na sedmo vprašanje odgovoriti, da je treba člen 5(5) Direktive 2001/29 razlagati tako, da če začasna dejanja reproduciranja, opravljena med procesom zbiranja podatkov, kot so ta v postopku v glavni stvari, izpolnjujejo vse pogoje iz člena 5(1) te direktive, je treba šteti, da izpolnjujejo pogoj, v skladu s katerim dejanja reproduciranja ne smejo biti v nasprotju z običajno uporabo dela in tudi ne smejo nerazumno posegati v zakonite interese imetnika pravic.
Stroški
Ker je ta postopek za stranke v postopku v glavni stvari ena od stopenj v postopku pred predložitvenim sodiščem, to odloči o stroških. Stroški, priglašeni za predložitev stališč Sodišču, ki niso stroški omenjenih strank, se ne povrnejo.
Iz teh razlogov je Sodišče (tretji senat) razsodilo:
Člen 5(1) Direktive 2001/29/ES Evropskega parlamenta in Sveta z dne 22. maja 2001 o usklajevanju določenih vidikov avtorske in sorodnih pravic v informacijski družbi je treba razlagati tako, da začasna dejanja reproduciranja, opravljena med procesom, imenovanim zbiranje podatkov“, kot so ta v postopku v glavni stvari,
izpolnjujejo pogoj, v skladu s katerim morajo biti ta dejanja sestavni in bistveni del tehnološkega procesa, ne glede na to, da pomenijo začetek in konec tega procesa ter zahtevajo človeško posredovanje;
so skladna s pogojem, v skladu s katerim morajo imeti dejanja reproduciranja samo en namen, in sicer zakonito uporabo zaščitenega dela ali predmeta sorodnih pravic;
izpolnjujejo pogoj, v skladu s katerim ta dejanja ne smejo imeti neodvisnega ekonomskega pomena, če izvedba teh dejanj ne omogoča ustvarjanja dodatnega dobička, ki presega dobiček v zvezi z zakonito uporabo zaščitenega dela, in če začasna dejanja reproduciranja ne privedejo do spremembe tega dela.
Člen 5(5) Direktive 2001/29 je treba razlagati tako, da če začasna dejanja reproduciranja, opravljena med procesom, imenovanim zbiranje podatkov“, kot so ta v postopku v glavni stvari, izpolnjujejo vse pogoje iz člena 5(1) te direktive, je treba šteti, da izpolnjujejo pogoj, v skladu s katerim dejanja reproduciranja ne smejo biti v nasprotju z običajno uporabo dela in tudi ne smejo nerazumno posegati v zakonite interese imetnika pravic.
Podpisi
DOMSTOLENS DOM (stora avdelningen)
den 24 januari 2012 ( *1 )
Socialpolitik — Direktiv 2003/88/EG — Artikel 7 — Rätt till årlig betald semester — Villkor för rätten föreskrivs i nationella bestämmelser — Arbetstagarens frånvaro — Ledighetens längd är beroende av frånvarons art — Nationella bestämmelser som strider mot direktiv 2003/88 — Den nationella domstolens roll”
I mål C-282/10,
angående en begäran om förhandsavgörande enligt artikel 267 FEUF, framställd av Cour de cassation (Frankrike) genom beslut av den 2 juni 2010, som inkom till domstolen den 7 juni 2010, i målet
Maribel Dominguez
mot
Centre informatique du Centre Ouest Atlantique,
Préfet de la région Centre,
meddelar
DOMSTOLEN (stora avdelningen)
sammansatt av ordföranden V. Skouris, avdelningsordförandena A. Tizzano, J.N. Cunha Rodrigues, K. Lenaerts och U. Lõhmus samt domarna A. Rosas, E. Levits (referent), A. Ó Caoimh, L. Bay Larsen, T. von Danwitz och A. Arabadjiev,
generaladvokat: V. Trstenjak,
justitiesekreterare: handläggaren R. Şereş,
efter det skriftliga förfarandet och förhandlingen den 17 maj 2011,
med beaktande av de yttranden som avgetts av:
Maribel Dominguez, genom H. Masse-Dessen och V. Lokiec, avocats,
Centre informatique du Centre Ouest Atlantique, genom D. Célice, avocat,
Frankrikes regering, genom G. de Bergues, A. Czubinski och N. Rouam, samtliga i egenskap av ombud,
Danmarks regering, genom S. Juul Jørgensen, i egenskap av ombud,
Nederländernas regering, genom C. Wissels och M. Noort, båda i egenskap av ombud,
Europeiska kommissionen, genom M. van Beek och M. Van Hoof, båda i egenskap av ombud,
och efter att den 8 september 2011 ha hört generaladvokatens förslag till avgörande,
följande
Dom
Begäran om förhandsavgörande avser tolkningen av artikel 7 i Europaparlamentets och rådets direktiv 2003/88/EG av den 4 november 2003 om arbetstidens förläggning i vissa avseenden (EUT L 299, s. 9).
Begäran har framställts i ett mål mellan Maribel Dominguez och hennes arbetsgivare, Centre informatique du Centre Ouest Atlantique (nedan kallat CICOA). Målet gäller Maribel Dominguez begäran att beviljas årlig betald semester som hon inte tagit ut under perioden mellan november 2005 och januari 2007 på grund av sjukskrivning till följd av en olycka, och i andra hand ett yrkande om kompensationsersättning.
Tillämpliga bestämmelser
Unionslagstiftningen
I artikel 1 i direktiv 2003/88 föreskrivs följande:
Ändamål och räckvidd
I detta direktiv föreskrivs minimikrav på säkerhet och hälsa vid förläggningen av arbetstiden.
Detta direktiv är tillämpligt på
minimitider för … årlig semester, …
...”
Artikel 7 i direktivet har följande lydelse:
Årlig semester
Medlemsstaterna skall vidta de åtgärder som behövs för att se till att varje arbetstagare får en årlig betald semester om minst fyra veckor i enlighet med vad som föreskrivs genom nationell lagstiftning eller praxis angående rätten till och beviljandet av en sådan semester.
Den årliga semestern får inte utbytas mot kontant ersättning, utom då anställningen avslutas.”
I artikel 15 i direktivet föreskrivs följande:
Gynnsammare bestämmelser
Detta direktiv skall inte påverka medlemsstaternas rätt att tillämpa eller införa lagar eller andra författningar som bättre skyddar arbetstagarnas hälsa och säkerhet eller underlättar eller tillåter tillämpningen av kollektivavtal eller avtal mellan arbetsmarknadens parter som bättre skyddar arbetstagarnas hälsa och säkerhet.”
I artikel 17 i direktiv 2003/88 föreskrivs att medlemsstaterna får göra avvikelser från vissa bestämmelser i direktivet. Avvikelser från artikel 7 i direktivet är inte tillåtna.
Den nationella lagstiftningen
I artikel L. 223-2, första stycket i lagen om arbete föreskrivs följande:
En arbetstagare, som under intjänandeåret kan styrka att vederbörande har varit anställd hos samma arbetsgivare under en tid som motsvarar minst en månads faktiskt arbete, har rätt till semester vars längd ska fastställas till två och en halv arbetsdagar per arbetsmånad, dock utan att det totala antalet semesterdagar får överstiga 30 arbetsdagar.”
Enligt artikel L. 223-4 i samma lag gäller följande:
Perioder som motsvarar fyra veckor eller 24 arbetsdagar ska likställas med en månads faktiskt arbete vid fastställandet av semesterns längd. Betalda semesterperioder, kompensationsledighet …, ledighet för kvinnor som har fött barn …, lediga dagar som har erhållits med anledning av arbetstidsförkortning och perioder som är begränsade till en sammanhängande tid på ett år då fullgörandet av anställningsavtalet är vilande på grund av ett olycksfall i arbetet eller yrkessjukdom ska anses utgöra perioder av faktiskt arbete. …”
I artikel XIV fjärde stycket i de standardföreskrifter som har bifogats det nationella kollektivavtalet för personal vid socialförsäkringsorgan föreskrivs följande:
Rätt till årlig semester föreligger inte under ett visst år vid frånvaro på grund av sjukdom eller långvarig sjukdom, som har föranlett ett uppehåll i arbetet som uppgår till eller överstiger tolv månader i följd, … Rätt till årlig semester uppstår på nytt när arbetet återupptas, varvid semesterns längd ska fastställas i proportion till den faktiska arbetstid som ännu inte har gett rätt till årlig semester.”
Målet vid den nationella domstolen och tolkningsfrågorna
Maribel Dominguez är sedan år 1987 anställd av CICOA och omfattas av det nationella kollektivavtalet för personal vid socialförsäkringsorgan. Efter att Maribel Dominguez hade råkat ut för en olycka på vägen från bostaden till arbetsplatsen var hon sjukskriven mellan den 3 november 2005 och den 7 januari 2007.
Maribel Dominguez väckte talan vid arbetsdomstol och överklagade därefter till Cour d’appel de Limoges för att beviljas 22,5 dagars betald semester för denna period och i andra hand utbetalning av en kompensationsersättning.
Sedan båda domstolarna ogillat hennes talan överklagade Maribel Dominguez till Cour de cassation. Hon har gjort gällande att olyckan på vägen till arbetet är ett olycksfall i arbetet som omfattas av samma regler som den sistnämnda olyckstypen. Med tillämpning av artikel L. 223-4 i lagen om arbete ska den period då hennes anställningsavtal var vilande på grund av olyckan på vägen till arbetet således jämställas med faktisk arbetstid vid beräkningen av betald ledighet.
Mot bakgrund av domstolens praxis avseende artikel 7 i direktiv 2003/88 hyser Cour de cassation tvivel angående huruvida de relevanta nationella bestämmelserna är förenliga med nämnda artikel.
Cour de cassation beslutade under dessa förhållanden att vilandeförklara målet och hänskjuta följande tolkningsfrågor till domstolen:
1)
Ska artikel 7.1 i direktiv 2003/88 … tolkas så, att den utgör hinder för nationella bestämmelser eller nationell praxis som innebär att det som villkor för rätten till årlig betald semester krävs att det utförs faktiskt arbete under minst tio dagar (eller en månad) under intjänandeperioden?
Om fråga 1 ska besvaras jakande: Är den nationella domstolen enligt artikel 7 i direktiv 2003/88 … – vilken medför en särskild skyldighet för arbetsgivaren, genom att den ger en arbetstagare som av hälsoskäl är frånvarande under en tid som uppgår till eller överstiger ett år rätt till betald semester – skyldig att, i en tvist mellan enskilda, underlåta att tillämpa en oförenlig nationell bestämmelse som i det fallet innebär att det, som villkor för rätten till årlig betald semester krävs, att faktiskt arbete har utförts under minst tio dagar under intjänandeåret?
Har arbetstagarna, eftersom det i artikel 7 i direktiv 2003/88… inte görs någon åtskillnad mellan arbetstagarna beroende på om deras frånvaro från arbetet under intjänandeperioden har orsakats av ett olycksfall i arbetet, en yrkessjukdom, ett olycksfall på väg till eller från arbetet eller en sjukdom som inte är yrkesrelaterad, enligt denna artikel rätt till betald semester som är lika lång oavsett orsaken till deras frånvaro av hälsoskäl, eller ska denna artikel tolkas så, att den inte utgör hinder för att längden på den betalda semestern kan variera beroende på orsaken till arbetstagarens frånvaro, eftersom det i den nationella lagen under vissa villkor föreskrivs en längd på den årliga betalda semestern som överstiger den minimilängd på fyra veckor som föreskrivs i direktiv [2003/88]?”
Prövning av den första frågan
Den nationella domstolen har ställt den första frågan för att få klarhet i huruvida artikel 7.1 i direktiv 2003/88 ska tolkas så, att den utgör hinder för nationella bestämmelser eller nationell praxis, som innebär att rätten till årlig betald semester är underställd villkoret att det utförs faktiskt arbete under minst tio dagar eller en månad under intjänandeperioden.
Det följer av fast rättspraxis att varje arbetstagares rätt till årlig betald semester måste betraktas som en princip av särskild betydelse i unionens sociala regelverk. Undantag från denna princip får därför inte göras, och de behöriga nationella myndigheternas genomförande av denna princip får endast ske inom de gränser som uttryckligen uppställs i rådets direktiv 93/104/EG av den 23 november 1993 om arbetstidens förläggning i vissa avseenden (EGT L 307, s. 18), kodifierat genom direktiv 2003/88 (se dom av den 26 juni 2001 i mål C-173/99, BECTU, REG 2001, s. I-4881, punkt 43, av den 20 januari 2009 i de förenade målen C-350/06 och C-520/06, Schultz-Hoff m.fl., REG 2009, s. I-179, punkt 22, och av den 22 november 2011 i mål C-214/10, KHS, ännu ej publicerat i rättsfallssamlingen, punkt 23).
Direktiv 93/104 ska följaktligen tolkas så, att det utgör hinder för att medlemsstaterna ensidigt begränsar den rätt till årlig betald semester som alla arbetstagare har genom att tillämpa ett villkor för den nämnda rättigheten som leder till att vissa arbetstagare utestängs från rättigheten (domen i det ovannämnda målet BECTU, punkt 52).
Medlemsstaterna får förvisso i sin interna lagstiftning fastställa villkoren för hur rätten till årlig betald semester ska utövas och genomföras. Det får dock inte uppställas något som helst villkor för själva uppkomsten av denna rättighet (domen i det ovannämnda målet Schultz-Hoff m.fl., punkt 46).
De verkställighets- och tillämpningsföreskrifter som är nödvändiga för att genomföra bestämmelserna i direktiv 93/104, vilket kodifierades genom direktiv 2003/88, kan således innehålla vissa skillnader vad gäller villkoren för utövande av rätten till årlig betald semester Enligt detta direktiv är det emellertid inte tillåtet för medlemsstaterna att utestänga någon från själva uppkomsten av en rätt som uttryckligen har tillerkänts alla arbetstagare (domarna i de ovannämnda målen BECTU, punkt 55, och Schultz-Hoff m.fl., punkt 47).
I direktiv 2003/88 görs dessutom inte någon åtskillnad mellan arbetstagare som är frånvarande från arbetet på grund av sjukledighet under intjänandeperioden och de som verkligen har arbetat under denna period (se domen i det ovannämnda målet Schultz-Hoff m.fl., punkt 40). Av detta följer att när det gäller arbetstagare som är sjukskrivna i vederbörlig ordning kan en medlemsstat inte som villkor för den rätt till årlig betald semester som enligt direktivet tillkommer alla arbetstagare föreskriva att arbetstagarna faktiskt måste ha arbetat under den intjänandeperiod som fastställts av nämnda stat (domen i det ovannämnda målet Schultz-Hoff m.fl., punkt 41).
Av vad som anförts ovan följer att artikel 7.1 i direktiv 2003/88 ska tolkas så, att den utgör hinder för nationella bestämmelser eller nationell praxis, som innebär att rätten till årlig betald semester är underställd villkoret att faktiskt arbete har utförts under en period om minst tio dagar eller en månad under intjänandeperioden.
Prövning av den andra frågan
Den hänskjutande domstolen har ställt den andra frågan för att få klarhet i huruvida artikel 7 i direktiv 2003/88 ska tolkas så, att en nationell bestämmelse som uppställer som villkor för rätten till årlig betald semester att en minimiperiod av faktiskt arbete har utförts under intjänandeperioden, i strid med nämnda artikel 7, inte ska tillämpas i en tvist mellan enskilda.
Domstolen erinrar inledningsvis om att frågan huruvida en nationell bestämmelse, för det fall den strider mot unionsrätten, inte ska tillämpas endast uppstår om det inte är möjligt att tolka bestämmelsen på ett sätt som är förenligt med unionsrätten.
Av fast rättspraxis framgår att de nationella domstolarna vid tillämpningen av nationell rätt är skyldiga att i den utsträckning det är möjligt tolka denna mot bakgrund av direktivets ordalydelse och syfte så att det resultat som avses i direktivet uppnås och, därmed, följa artikel 288 tredje stycket FEUF. Denna skyldighet att göra en direktivkonform tolkning av nationell rätt följer av EUF-fördragets systematik, eftersom den gör det möjligt för de nationella domstolarna att inom ramen för sin behörighet säkerställa att unionsrätten ges full verkan när de avgör tvister som anhängiggjorts vid dem (se, bland annat, dom av den 5 oktober 2004 i de förenade målen C-397/01-C-403/01, Pfeiffer m.fl., REG 2004, s. I-8835, punkt 114, av den 23 april 2009 i de förenade målen C-378/07-C-380/07, Angelidaki m.fl., REG 2009, s. I-3071, punkterna 197 och 198, samt domen av den 19 januari 2010 i mål C-555/07, Kücükdeveci, REU 2010, s. I-365, punkt 48).
Principen om direktivkonform tolkning av nationell rätt har förvisso vissa begränsningar. Den nationella domstolens skyldighet att beakta ett direktivs innehåll vid tolkningen och tillämpningen av relevanta bestämmelser i nationell rätt begränsas således av allmänna rättsprinciper och den kan inte tjäna som grund för att nationell rätt tolkas contra legem (se dom av den 15 april 2008 i mål C-268/06, Impact, REG 2008, s. I-2483, punkt 100, samt domen i det ovannämnda målet Angelidaki m.fl., punkt 199).
Den hänskjutande domstolen anser att den står inför en sådan begränsning i det nationella målet. Enligt nämnda domstol kan artikel L. 223-2, första stycket i lagen om arbete, enligt vilken rätten till årlig betald semester är underställd ett krav på att minst en månads faktiskt arbete har utförts under beräkningsperioden, inte tolkas på ett sätt som är förenligt med artikel 7 i direktiv 2003/88.
Principen om direktivkonform tolkning innebär icke desto mindre att de nationella domstolarna ska göra allt som ligger inom deras behörighet, med hänsyn till den nationella rätten i sin helhet och med tillämpning av de tolkningsmetoder som är erkända i nationell rätt, för att säkerställa att det aktuella direktivet ges full verkan och för att uppnå ett resultat som är förenligt med direktivets syfte (se dom av den 4 juli 2006 i mål C-212/04, Adeneler m.fl., REG 2006, s. I-6057, punkt 111, samt domen i det ovannämnda målet Angelidaki m.fl., punkt 200).
I det nationella målet utgör artikel L. 223-4 i lagen om arbete – enligt vilken vissa typer av frånvaro från arbetet anses berättiga till undantag från kravet på att faktiskt arbete ska ha utförts under intjänandeperioden – en väsentlig del av den nationella rätten som de nationella domstolarna ska beakta.
Om den hänskjutande domstolen, för att ge artikel 7 i direktiv 2003/88 full verkan, skulle tolka artikel L. 223-4 i lagen om arbete så att en frånvaroperiod på grund av en olycka på vägen till arbetet ska likställas med en frånvaroperiod på grund av olycksfall i arbetet, skulle nämnda domstol inte ställas inför den begränsning som följer av en direktivkonform tolkning av artikel L. 223-2 i lagen om arbete, som nämns ovan i punkt 26.
Det ska i detta avseende preciseras att artikel 7 i direktiv 2003/88 inte gör någon åtskillnad mellan de arbetstagare som är frånvarande under intjänandeperioden på grund av sjukskrivning och dem som verkligen har arbetat under denna period (se punkt 20 i denna dom). Detta innebär att en medlemsstat inte kan underställa rätten till årlig betald semester – för en arbetstagare som under intjänandeperioden har varit frånvarande från arbetet av hälsoskäl – ett krav på att vederbörande ska ha utfört faktiskt arbete under denna period. Enligt artikel 7 i direktiv 2003/88 kan således inte någon arbetstagares rätt till årlig betald semester om minst fyra veckor påverkas, oavsett om vederbörande har varit sjukledig under intjänandeperioden på grund av ett olycksfall på arbetsplatsen eller någon annanstans eller till följd av sjukdom, oavsett slag eller orsak.
Av det ovan anförda följer att det ankommer på den hänskjutande domstolen att kontrollera om den – med beaktande av den nationella rätten i dess helhet, i synnerhet artikel L. 223-4 i lagen om arbete, och med tillämpning av de tolkningsmetoder som erkänns i nationell rätt –, för att säkerställa att direktiv 2003/88 ges full verkan och för att uppnå ett resultat som är förenligt med direktivets syfte, kan tolka nationell rätt på ett sätt som gör det möjligt att likställa en arbetstagares frånvaro på grund av en olycka som inträffat på vägen till arbetet med en av de frånvarotyper som nämns i artikel L. 223-4 i lagen om arbete.
Om en sådan tolkning inte är möjlig, ska det prövas om artikel 7.1 i direktiv 2003/88 har direkt effekt och, om så är fallet, om Maribel Dominguez kan åberopa denna gentemot svarandena i det nationella målet, i synnerhet hennes arbetsgivare CICOA, med hänsyn till deras rättsliga natur.
Det följer härvid av domstolens fasta praxis att enskilda, i alla de fall då bestämmelserna i ett direktiv med avseende på innehållet framstår som ovillkorliga och tillräckligt precisa, har rätt att åberopa dem inför den nationella domstolen gentemot staten, när denna inte har införlivat direktivet med nationell rätt inom fristen eller inte har införlivat direktivet på ett korrekt sätt (se, bland annat, domen i det förenade målet Pfeiffer m.fl., punkt 103 och där angiven rättspraxis).
Artikel 7 i direktiv 2003/88 uppfyller emellertid dessa kriterier, eftersom medlemsstaterna i otvetydiga ordalag åläggs en skyldighet som ska leda till ett preciserat resultat och som inte är förenad med något villkor angående tillämpningen av den regel som föreskrivs däri, nämligen att ge alla arbetstagare rätt till en årlig betald semester om minst fyra veckor.
Även om artikel 7 i direktiv 2003/88 ger medlemsstaterna ett visst utrymme för skönsmässig bedömning när de fastställer villkoren för att erhålla och beviljas den rätt till årlig betald semester som föreskrivs i direktivet, påverkar dessa omständigheter inte den precisa och ovillkorliga karaktären som kännetecknar den skyldighet som föreskrivs i artikeln. Det ska noteras att artikel 7 i direktiv 2003/88 inte ingår bland de bestämmelser i direktivet som det enligt artikel 17 är möjligt att avvika från. Det är således möjligt att fastställa det minimiskydd som medlemsstaterna under alla omständigheter ska genomföra enligt artikel 7 (se, analogt, domen i det ovannämnda målet Pfeiffer m.fl., punkt 105).
Eftersom artikel 7.1 i direktiv 2003/88 uppfyller villkoren för att ha direkt effekt, konstaterar domstolen dessutom att CICOA, en av svarandena i det nationella målet, som är Maribel Dominguez arbetsgivare, är ett socialförsäkringsorgan.
Det är förvisso riktigt att ett direktiv enligt fast rättspraxis inte i sig kan medföra skyldigheter för en enskild och det kan således inte som sådant åberopas gentemot denne (se, bland annat, dom av den 14 juli 1994 i mål C-91/92, Faccini Dori, REG 1994, s. I-3325, punkt 20, svensk specialutgåva, volym 16, s. I-1, av den 7 mars 1996 i mål C-192/94, El Corte Inglés, REG 1996, s. I-1281, punkt 15, domarna i de ovannämnda målen Pfeiffer m.fl., punkt 108, och Kücükdeveci, C-555/07, REU 2010, s. I-365, punkt 46).
Det ska emellertid påpekas att när enskilda rättssubjekt har möjlighet att stödja sig på ett direktiv, vid talan inte mot en enskild utan mot staten, kan de dessutom göra detta oavsett om staten agerar i egenskap av arbetsgivare eller myndighet. I båda fallen är det nämligen angeläget att staten hindras från att dra nytta av sin underlåtenhet att följa unionsrätten (se, bland annat, dom av den 26 februari 1986 i mål C-152/84, Marshall, REG 1986, s. 723, punkt 49, svensk specialutgåva, volym 8, s. 457, av den 12 juli 1990 i mål C-188/89, Foster m.fl., REG 1990, s. I-3313, punkt 17, svensk specialutgåva, volym 10, s. 479, samt av den 14 september 2000 i mål C-343/98, Collino och Chiappero, REG 2000, s. I-6659, punkt 22).
Bland de organ gentemot vilka sådana bestämmelser i ett direktiv som kan ha direkt effekt kan åberopas ingår ett organ som, oavsett sin rättsliga form, i enlighet med en av staten antagen rättsakt har fått i uppdrag att utöva offentlig serviceverksamhet under statens tillsyn och som med anledning härav har särskilda befogenheter utöver dem som följer av de rättsregler som gäller i förhållandet mellan enskilda (se, bland annat, domarna i de ovannämnda målen Foster m.fl., punkt 20, Collino och Chiappero, punkt 23, och dom av den 19 april 2007 i mål C-356/05, Farrell, REG 2007, s. I-3067, punkt 40).
Det ankommer således på den nationella domstolen att kontrollera om artikel 7.1 i direktiv 2003/88 kan åberopas gentemot CICOA.
Om så är fallet innebär artikel 7 i direktiv 2003/88, som uppfyller villkoren för att ha direkt effekt, att den nationella domstolen ska underlåta att tillämpa alla nationella bestämmelser som strider mot den.
Om så inte skulle vara fallet erinrar domstolen om att även om en direktivsbestämmelse som syftar till att tillerkänna enskilda rättigheter eller ålägga dem skyldigheter är klar, precis och ovillkorlig kan den inte som sådan tillämpas inom ramen för en tvist som enbart rör enskilda (se domen i det ovannämnda målet Pfeiffer m.fl., punkt 109).
I en sådan situation kan den part som lidit skada till följd av att nationell rätt inte är förenlig med unionsrätten dock åberopa rättspraxis i domen av den 19 november 1991 i de förenade målen C-6/90 och C-9/90, Francovich m.fl. (REG 1991, s. I-5357; svensk specialutgåva, volym 11, s. 435) för att i förekommande fall erhålla ersättning för den lidna skadan.
Den andra frågan ska följaktligen besvaras enligt följande:
Det ankommer på den hänskjutande domstolen att kontrollera om den – för att säkerställa att artikel 7 i direktiv 2003/88 ges full verkan och för att uppnå ett resultat som är förenligt med direktivets syfte – kan tolka nationell rätt på ett sätt som gör det möjligt att likställa en arbetstagares frånvaro på grund av en olycka som inträffat på vägen till arbetet med en av de frånvarotyper som nämns i artikel L. 223-4 i lagen om arbete. Detta ska ske med beaktande av nationell rätt i dess helhet, i synnerhet nämnda artikel L. 223-4, och med tillämpning av de tolkningsmetoder som erkänns i nationell rätt.
Om en sådan tolkning inte är möjlig ankommer det på den nationella domstolen att, med hänsyn till den rättsliga naturen hos svarandena i det nationella målet, kontrollera om den direkta effekten av artikel 7.1 i direktiv 2003/88 kan åberopas mot dem.
Om den nationella domstolen inte kan uppnå det resultat som föreskrivs i artikel 7 i direktiv 2003/88, kan den part som lidit skada till följd av att nationell rätt inte är förenlig med unionsrätten dock åberopa domen i målet Francovich m.fl., för att i förekommande fall erhålla ersättning för den lidna skadan.
Den tredje frågan
Den hänskjutande domstolen har ställt den tredje frågan för att få klarhet i huruvida artikel 7 i direktiv 2003/88 ska tolkas så, att den utgör hinder för en nationell bestämmelse vari det föreskrivs, beroende på orsaken till arbetstagarens sjukfrånvaro, en årlig betald semester som överstiger eller är lika med den minimilängd på fyra veckor som garanteras i direktivet.
Domstolen erinrar härvid, i likhet med vad som konstateras i punkt 30 i denna dom, om att det i artikel 7 i direktiv 2003/88 inte görs någon åtskillnad utifrån orsaken till att en arbetstagare är frånvarande på grund av en sjukskrivning som skett i vederbörlig ordning. Alla arbetstagare har nämligen rätt till en årlig betald semester om minst fyra veckor, oavsett om arbetstagaren sjukskrivits till följd av ett olycksfall på arbetsplatsen eller någon annanstans eller till följd av sjukdom, oavsett slag eller orsak.
Vad som konstaterades i föregående punkt innebär emellertid inte att direktiv 2003/88 utgör hinder för nationella bestämmelser vari föreskrivs en rätt till årlig betald semester under mer än fyra veckor som beviljas och erhålles enligt villkor som fastställs i nationell rätt. Detta påpekade såväl generaladvokaten i punkt 178 i sitt förslag till avgörande som Europeiska kommissionen i sin skriftliga inlaga.
Det följer nämligen uttryckligen av ordalydelsen i artiklarna 1.1, 1.2 a, 7.1 och 15 i direktiv 2003/88 att ändamålet med direktivet endast är att föreskriva minimikrav på säkerhet och hälsa vid förläggningen av arbetstiden och att direktivet inte påverkar medlemsstaternas rätt att tillämpa nationella bestämmelser som bättre skyddar arbetstagarna.
Det är således tillåtet för medlemsstaterna att föreskriva att rätten till årlig betald semester enligt nationell rätt ska variera beroende på orsaken till att arbetstagaren är frånvarande av hälsoskäl, under förutsättning att den alltid överstiger eller är lika med den minimilängd på fyra veckor som föreskrivs i artikel 7 i direktivet.
Det följer av vad som anförts att artikel 7.1 i direktiv 2003/88 ska tolkas så, att den inte utgör hinder för en nationell bestämmelse vari det föreskrivs, beroende på orsaken till arbetstagarens sjukfrånvaro, en årlig betald semester som överstiger eller är lika med den minimilängd på fyra veckor som garanteras i direktivet.
Rättegångskostnader
Eftersom förfarandet i förhållande till parterna i målet vid den nationella domstolen utgör ett led i beredningen av samma mål, ankommer det på den nationella domstolen att besluta om rättegångskostnaderna. De kostnader för att avge yttrande till domstolen som andra än nämnda parter har haft är inte ersättningsgilla.
Mot denna bakgrund beslutar domstolen (stora avdelningen) följande:
Artikel 7.1 i Europaparlamentets och rådets direktiv 2003/88/EG av den 4 november 2003 om arbetstidens förläggning i vissa avseenden ska tolkas så, att den utgör hinder för nationella bestämmelser eller nationell praxis, som innebär att rätten till årlig betald semester är underställd villkoret att faktiskt arbete har utförts under en period om minst tio dagar eller en månad under intjänandeperioden.
Det ankommer på den hänskjutande domstolen att kontrollera om den – för att säkerställa att artikel 7 i direktiv 2003/88 ges full verkan och för att uppnå ett resultat som är förenligt med direktivets syfte – kan tolka nationell rätt på ett sätt som gör det möjligt att likställa en arbetstagares frånvaro på grund av en olycka som inträffat på vägen till arbetet med en av de frånvarotyper som nämns i artikel L. 223-4 i lagen om arbete. Detta ska ske med beaktande av nationell rätt i dess helhet, i synnerhet nämnda artikel L. 223-4, och med tillämpning av de tolkningsmetoder som erkänns i nationell rätt.
Om en sådan tolkning inte är möjlig ankommer det på den nationella domstolen att, med hänsyn till den rättsliga naturen hos svarandena i det nationella målet, kontrollera om den direkta effekten av artikel 7.1 i direktiv 2003/88 kan åberopas mot dem.
Om den nationella domstolen inte kan uppnå det resultat som föreskrivs i artikel 7 i direktiv 2003/88, kan den part som lidit skada till följd av att nationell rätt inte är förenlig med unionsrätten dock åberopa rättspraxis i domen av den 19 november 1991 i de förenade målen C-6/90 och C-9/90, Francovich m.fl., för att i förekommande fall erhålla ersättning för den lidna skadan.
Artikel 7.1 i direktiv 2003/88 ska tolkas så, att den inte utgör hinder för en nationell bestämmelse vari det föreskrivs, beroende på orsaken till arbetstagarens sjukfrånvaro, en årlig betald semesterperiod som överstiger eller är lika med den minimilängd på fyra veckor som garanteras i direktivet.
Underskrifter
DOMSTOLENS DOM (första avdelningen)
den 2 februari 2012 ( *1 )
Konventionen med stadga för Europaskolorna — Tolkning och tillämpning av artiklarna 12.4 a och 25.1 — Rätt för de utstationerade lärarna att få tillträde till samma karriär- och löneutvecklingsmöjligheter som deras nationella motsvarigheter — Vissa lärare som har utstationerats av Förenade kungariket vid Europaskolorna är uteslutna från tillträde till mer fördelaktiga löneskalor och andra tilläggsbetalningar som erbjuds deras nationella motsvarigheter — Oförenlighet med artiklarna 12.4 a och 25.1”
I mål C-545/09,
angående en talan enligt artikel 26 i konventionen med stadga för Europaskolorna, väckt den 22 december 2009,
Europeiska kommissionen, företrädd av J. Currall och B. Eggers, båda i egenskap av ombud, med delgivningsadress i Luxemburg,
sökande,
mot
Förenade konungariket Storbritannien och Nordirland, företrätt av H. Walker, i egenskap av ombud, och J. Coppel, barrister,
svarande,
meddelar
DOMSTOLEN (första avdelningen)
sammansatt av avdelningsordföranden A. Tizzano samt domarna A. Borg Barthet, M. Ilešič (referent), J.-J. Kasel och M. Berger,
generaladvokat: P. Mengozzi,
justitiesekreterare: handläggaren K. Sztranc-Sławiczek,
efter det skriftliga förfarandet och förhandlingen den 4 maj 2011,
och efter att den 7 juli 2011 ha hört generaladvokatens förslag till avgörande,
följande
Dom
Europeiska kommissionen har yrkat att domstolen ska fastställa att artikel 12.4 a i konventionen med stadga för Europaskolorna av den 21 juni 1994 (EGT L 212, s. 3) (nedan kallad konventionen) ska tolkas och tillämpas så, att den garanterar att lärare som har utstationerats av en medlemsstat, under den tid som utstationeringen varar, får tillträde till samma karriär- och löneutvecklingsmöjligheter som lärare som tjänstgör inom den medlemsstatens territorium samt att det är oförenligt med artiklarna 12.4 a och 25.1 i konventionen att utesluta vissa lärare som har utstationerats av Förenade konungariket Storbritannien och Nordirland, under den tid som utstationeringen varar, från det tillträde, som lärare anställda vid offentliga skolor i England och Wales har, till mer fördelaktiga löneskalor (bland annat ”threshold pay”, ”excellent teacher system” och ”advanced skills teachers”) och andra tilläggsbetalningar (som ”teaching and learning responsibility payments”) samt uppflyttning inom den befintliga löneskalan.
Tillämpliga bestämmelser
Konventionen och stadgan för den utstationerade personalen
Europaskolorna inrättades ursprungligen med stöd av två rättsakter, dels stadgan för Europaskolan, som undertecknades i Luxemburg den 12 april 1957 (Recueil des traités des Nations unies, volym 443, s. 129), dels protokollet om grundande av Europaskolor, vilket upprättats med hänvisning till nämnda stadga och som undertecknades i Luxemburg den 13 april 1962 (Recueil des traités des Nations unies, volym 752, s. 267).
Dessa rättsakter ersattes av den konvention som trädde i kraft den 1 oktober 2002 och som är den konvention som just nu äger tillämpning. Till skillnad från de ursprungliga rättsakterna, där endast medlemsstaterna var parter, ingicks konventionen även av Europeiska gemenskaperna, vilka bemyndigats härför genom rådets beslut 94/557/EG, Euratom av den 17 juni 1994 om bemyndigande för Europeiska gemenskapen och Europeiska atomenergigemenskapen att underteckna och sluta konventionen med stadga för Europaskolorna (EGT L 212, s. 1; svensk specialutgåva, område 16, volym 2, s. 81).
I det tredje skälet i konventionen anges följande:
som beaktar att Europaskolsystemet är en särskild typ av skolsystem och som beaktar att det utgör en form av samarbete mellan medlemsstaterna och mellan dem och Europeiska gemenskaperna och som samtidigt helt erkänner medlemsstaternas ansvar för undervisningens innehåll och organisationen av sina utbildningssystem, och för sin kulturella och språkliga mångfald”.
I artikel 3.2 i konventionen föreskrivs följande:
Undervisningen skall ske genom lärare som är utsända eller utnämnda av medlemsstaterna i enlighet med beslut som fattats av styrelsen enligt det förfarande som fastställs i artikel 12.4.”
I artikel 12.4 a i konventionen, som hör till avdelning II med rubriken ”Skolornas organ”, föreskrivs följande:
I administrativa frågor skall styrelsen ha följande uppgifter:
...
Den skall varje år på förslag av skolinspektörsnämnderna besluta om behovet av lärarpersonal genom inrättande eller indragning av tjänster. Den skall säkerställa en rättvis fördelning av tjänster bland medlemsstaterna. Den skall med regeringarna lösa frågor angående utnämning eller utstationering av lärare på de olika nivåerna och studievägledare i skolan. Personalen skall behålla de rättigheter ifråga om befordring och pension som garanteras enligt nationella regler.”
I artikel 25 i konventionen föreskrivs följande:
Skolornas budget skall finansieras genom
bidrag från medlemsstaterna genom fortsatt utbetalning av lön till utsända eller utnämnda lärare och, vid behov, ett finansiellt bidrag som enhälligt beslutats av styrelsen,
bidrag från Europeiska gemenskaperna avsett att täcka skillnaden mellan den totala utgiftssumman för skolorna och summan av andra inkomster,
bidrag från icke-gemenskapsorganisationer med vilka styrelsen har slutit avtal,
skolans egen inkomst, dvs. skolavgifterna som debiteras föräldrarna av styrelsen,
diverse inkomster.
Reglerna för bidrag från Europeiska gemenskaperna skall fastställas i en särskild överenskommelse mellan styrelsen och kommissionen.”
Enligt artikel 26 i konventionen ska ”Europeiska gemenskapernas domstol … ensam ha behörighet i tvister mellan de fördragsslutande parterna, vad avser tolkning och tillämpning av denna konvention, vilka inte har lösts av styrelsen.”
På grundval av artikel 12.1 i konventionen antog styrelsen stadgan för den utstationerade personalen vid Europaskolorna (nedan kallad stadgan för den utstationerade personalen), vilken bland annat innehåller bestämmelser om lön och arbetsvillkor för lärare vid Europaskolorna.
Enligt artikel 10.1 i stadgan för den utstationerade personalen ska de utstationerade lärarna besitta de kvalifikationer och uppfylla de nödvändiga villkor som erfordras för att inneha motsvarande befattningar i de länder de kommer från. I artikel 30 första stycket, som återfinns i kapitel III i stadgan med rubriken ”Utvärdering”, föreskrivs följande. ”Personalmedlems sakkunskap, effektivitet och anpassning i tjänsten är för undervisnings- och övervakningspersonal liksom för biträdande rektorer föremål för en utvärderingsrapport, som skall upprättas i lika mån av rektor som av den nationella inspektören, enligt de bestämmelser som finns fastställda i tillämpningsbestämmelserna. Om meningsskiljaktighet skulle föreligga, skall den nationella inspektörens rapport ha företräde.”
Enligt artikel 49 i stadgan uppbär den utstationerade personalen de nationella löner som behöriga nationella myndigheter utbetalar samt ett tillägg motsvarande skillnaden mellan den lön som föreskrivs i stadgan och värdet av den nationella lönen med avdrag för obligatoriska sociala avgifter. Tillägget betalas ut av Europaskolan (nedan kallat det europeiska tillägget).
En personalmedlem som slutgiltigt lämnar sin tjänst har dessutom – förutsatt att detta inte sker till följd av en disciplinåtgärd – enligt artikel 72.1 i stadgan rätt till ett avgångsvederlag som står i proportion till den faktiska tjänstgöringstiden upp till den maximala perioden om nio år. Avgångsvederlaget beräknas enligt artikel 72.2 som antalet tjänstgöringsår multiplicerat med differensen mellan en och en halv månad med den sista europeiska grundlönen korrigerad med den för ursprungslandet fastställda koefficienten, och en och en halv månad med den sista nationella grundlönen.
Stadgan innehåller däremot inget pensionssystem för utstationerade lärare, vilka under utstationeringen fortsätter att betala avgifter till sina nationella pensionssystem.
Bestämmelser som är tillämpliga på lärare som är anställda i England och Wales
I Förenade kungariket är utbildningssystemet föremål för en decentraliserad behörighet fördelad på tre separata regioner: England och Wales (som tillsammans utgör en region i detta avseende), Nordirland och Skottland. Arbetsvillkoren skiljer sig mellan dessa tre regioner.
I den region som utgörs av England och Wales – den enda region som är i fråga i den aktuella tvisten – är de flesta lärarna anställda vid någon av de statsunderstödda skolorna (”maintained schools”). Lön och arbetsvillkor för dessa lärare fastställs genom beslut av behörig minister, närmare bestämt i ett dokument avseende lön och villkor för skollärare (”School Teachers Pay and Conditions Document”, nedan kallat STPCD), som är bindande för alla anställningsavtal som ingås av en statsunderstödd skola.
Ett visst antal lärare är inte anställda vid statsunderstödda skolor utan vid andra typer av skolor, till exempel fristående statliga skolor som stöds av sponsorer (”academies”), privatskolor, Europaskolan i Culham eller skolor som drivs av utländska regeringar. För dessa skolor är formerna och villkoren för arbetet enligt STPCD fakultativa.
Löneskalorna i 2009 års version av STPCD ser i huvudsak ut som följer.
För lärarna finns det en grundlöneskala indelad i sex löneklasser. Det huvudsakliga kriteriet för att flyttas upp till nästa klass är erfarenhet mätt i antal tjänsteår. Bortsett från undantagsfall med otillfredsställande resultat sker uppflyttning inom denna löneskala således automatiskt.
År 2000 gjordes en generell löneökning på tre procent i England och Wales. Samtidigt gjordes en löneökning på sju procent på grundval av ett nytt system kallat ”threshold pay”. En lärare måste uppfylla vissa krav för att omfattas av det nya systemet.
Enligt detta system kan engelska och walesiska lärare som har nått grundlöneskalans högsta löneklass ansöka om tillämpningen av en övre löneskala (”post-threshold pay scale”). En lärare som vill ansöka om detta måste uppfylla vissa yrkesmässiga normer, styrka sina kvalifikationer och begära att få sin kompetens bedömd. Utvärderingarna görs av rektorerna. De yrkesmässiga normer som lärarna ska uppfylla anges i dokumentet ”Yrkesmässiga normer för lärare” (”Professional Standards for Teachers”). När en lärare omfattas av den övre löneskalan (och blivit ”post-threshold teacher”) handlar det inte om automatisk uppflyttning, utan eventuell uppflyttning sker på grundval av slutsatserna från årliga utvärderingssamtal.
Dessutom kan statsunderstödda skolor enligt STPCD inrätta tjänster för ”utmärkta lärare” (”excellent teachers”) och ”lärare med särskilda färdigheter” (”advanced skills teachers”), för vilka det finns separata löneskalor, samt tjänster som ger rätt till tilläggsbetalningar för undervisnings- och lärandeansvar (”teaching and learning responsibility payments”). En lärare kan inte samtidigt inneha flera av dessa tjänster.
För att få delta i ”excellent teacher scheme” måste en lärare ha befunnit sig i minst två år på den högsta av de tre nivåerna i ”post-threshold pay scale” och visa prov på specifik yrkeskompetens enligt vad som anges i ”Professional Standards for Teachers”. En lärare kan emellertid endast begära en utvärdering, som görs av utomstående personer, för detta ändamål i samband med att han eller hon söker en ledig ”excellent teacher”-tjänst vid sin egen skola. En ”excellent teacher” ska vid sidan av sina ordinarie undervisningsuppgifter också hjälpa andra lärare att bli effektivare och att förbättra sin undervisningskvalitet.
För att kunna komma i fråga för en ”advanced skills teacher”-tjänst behöver en lärare inte nödvändigtvis redan ha fått tillträde till ”post-threshold pay scale”, men han eller hon måste uppfylla ”post-threshold teacher standards” och särskilt de yrkesmässiga normer som gäller specifikt för ”advanced skills teachers” enligt vad som anges i ”Professional Standards for Teachers”. Utvärderingarna i detta avseende görs av utomstående personer. Dessa tjänster innebär ytterligare åtaganden som utförs till gagn för lärare från andra skolor.
För ”teaching and learning responsibility payments” kan slutligen alla undervisande lärare komma i fråga utan att det finns något krav på att de ska ha fått tillträde till ”post-threshold pay scale”. Dessa tilläggsbetalningar ges till lärare som tar på sig ”ett varaktigt kompletterande ansvar inom ramen för [skolans] personalstruktur”. Tanken är att ge kompensation för ansvar bland annat i fråga om att hjälpa elever utanför klassrummet eller att spela en drivande roll när det gäller ämnes- eller läroplansutveckling.
Bestämmelser som är tillämpliga på lärare som är utnämnda eller utstationerade av England och Wales vid Europaskolorna
Förenade kungarikets tjänster vid Europaskolorna är öppna för alla lärare med tillräckliga kvalifikationer, oberoende av huruvida de vid tidpunkten för utnämningen eller utstationeringen är anställda av en statsunderstödd skola, en privatskola, en skola utanför landets gränser eller till och med ingen utbildningsinrättning alls.
De lärare som är utstationerade av Förenade kungariket vid Europaskolorna behåller inte sin avtalsmässiga relation till sin tidigare arbetsgivare, utan ingår i samband med utstationeringen ett nytt anställningsavtal med ”Department for Children, Schools and Families” (ministeriet för barndoms-, skol- och familjefrågor, nedan kallat utbildningsministeriet).
I det anställningsavtalet anges det, när det gäller engelska och walesiska lärare, att STPCD inte är tillämpligt på lärare vid Europaskolorna. Det slås emellertid fast att de nationella löner som varje månad betalas ut till de utstationerade lärarna ska fastställas i enlighet med löneskalorna i STPCD och att dessa lärare ska ha rätt till årliga löneökningar som förhandlas fram på nationell nivå och är tillämpliga i kraft av STPCD. Det anges också att inga andra tillägg till den nationella lönen ska betalas ut och att en utstationerad lärare inte har rätt att, så länge tjänstgöringen vid Europaskolorna varar, ansöka om uppflyttning till en högre löneskala, tilläggsbetalning eller en annan ställning enligt STPCD. Slutligen slås det fast i anställningsavtalet att tjänstgöring vid en Europaskola ger rätt till pension enligt pensionssystemet för engelska och walesiska lärare och att avgifterna till det systemet kommer att grunda sig uteslutande på den nationella lönen.
Förfarandet före talans väckande
Med anledning av ett stort antal klagomål från berörda lärare och flera frågor från Europaparlamentets ledamöter har kommissionen sedan år 2000 flera gånger vänt sig till Förenade kungarikets olika utbildningsministrar vid respektive tidpunkt och påpekat att det är oförenligt med konventionen att förvägra brittiska lärare utstationerade vid Europaskolorna möjligheten att få tillträde till den nya löneskalan. Varken en första skriftväxling under åren 2000 och 2001 eller en andra under 2007 erbjöd någon lösning på meningsskiljaktigheterna. Då begärde kommissionen att frågan skulle tas upp vid sammanträdet för Europaskolornas styrelse den 20–22 oktober 2008. Den 20 november 2008 hölls en videokonferens mellan företrädare för kommissionen och utbildningsministeriet, men inte heller denna kunde överbrygga oenigheten. Den 13 januari 2009 ingav kommissionen en sista begäran till styrelsen i syfte att finna en lösning på situationen och meddelade samtidigt att den, om inget resultat uppnåddes, ansåg sig tvungen att väcka talan vid domstolen.
Frågan om tolkningen av artiklarna 12.4 a och 25.1 i konventionen diskuterades vid styrelsesammanträdet den 20–21 januari 2009. Efter mötet konstaterade styrelsen att den ”inte hade lyckats slita tvisten och noterade att kommissionen hade för avsikt att vända sig till domstolen för att där väcka talan om tolkning och tillämpning mot Förenade kungariket med stöd av artikel 26 i konventionen i kombination med artiklarna 10 EG och 39 EG”.
Under dessa förhållanden beslutade kommissionen att väcka förevarande talan.
Talan
Kommissionen har yrkat att domstolen, med stöd av artikel 26 i konventionen, ska uttala sig om hur artikel 12.4 a sista meningen i konventionen ska tolkas samt pröva huruvida Förenade kungariket tillämpar den bestämmelsen korrekt, särskilt när det gäller lärare som har utstationerats av England och Wales vid Europaskolorna, och således uppfyller de förpliktelser som följer av den bestämmelsen och av artikel 25.1 i konventionen.
Tolkningen av artikel 12.4 a sista meningen i konventionen
Parternas argument
Kommissionen anser att sista meningen i artikel 12.4 a i konventionen ålägger medlemsstaterna en skyldighet att garantera att de utstationerade lärarna behåller de rättigheter i fråga om befordring och pension som garanteras enligt nationella regler. Denna konvention tilldelar, på grund av detta och i detta avseende, de utstationerade lärarna en rättighet.
Denna tolkning bekräftas enligt kommissionen av bestämmelsens klara och ovillkorliga lydelse samt av sammanhanget och bestämmelsens syfte, vilket är att lärarna inte ska missgynnas av sin utstationering.
Kommissionen har också gjort gällande att termen ”befordring” ska ges en fristående tolkning och avser att omfatta de olika nationella ersättningssystem som är tillämpliga på lärare vid utstationering. Termens stora räckvidd bekräftas av en analys av de olika språkversionerna.
Förenade kungariket anser däremot att artikel 12.4 a i konventionen riktar sig uteslutande till styrelsen och inte ålägger medlemsstaterna någon skyldighet.
Enligt Förenade kungariket bekräftas denna tolkning dels av bestämmelsens lydelse, som hör till avdelning II med rubriken ”Skolornas organ” i vilken ingen bestämmelse ålägger medlemsstaterna några skyldigheter, dels av den hänvisning som i artikel 3.2 i konventionen görs till artikel 12 i konventionen.
Enligt Förenade kungariket innebär artikel 12.4 a i konventionen att styrelsen vid utövandet av sina administrativa funktioner måste iaktta nationella regler i fråga om befordran och pension. Det skulle nämligen enligt Förenade kungariket inte vara rimligt att anse att konventionen ålägger medlemsstaterna att följa sin egen lagstiftning.
Enligt Förenade kungariket skulle det också strida mot artikel 165.1 FEUF, enligt vilken medlemsstaterna själva bestämmer hur deras utbildningssystem ska vara organiserade, om konventionen ålade medlemsstaterna en skyldighet att tillerkänna lärare som har utstationerats eller utnämnts vid Europaskolorna rättigheter som dessa lärare inte kan göra anspråk på enligt nationell lagstiftning.
Dessutom har denna medlemsstat gjort gällande att termen ”befordring”, i den betydelse som är allmänt vedertagen i Förenade kungariket, uteslutande avser att en lärare går vidare till en högre administrativ tjänst med större ansvar inom skolornas organisation, exempelvis en tjänst som rektor eller biträdande rektor (”head teacher” eller ”deputy head teacher”). När det gäller termerna ”rättigheter som garanteras” enligt nationella regler, har Förenade kungariket i huvudsak hävdat att dessa termer ska tolkas bokstavligt och restriktivt. En befordring – som inte automatiskt följer av tjänstetid utan som läraren måste ansöka om och som läraren åtnjuter endast om han eller hon uppfyller vissa krav – utgör således inte en rättighet som garanteras enligt nationella regler.
Domstolens bedömning
Meningsskiljaktigheterna mellan kommissionen och Förenade kungariket avseende tolkningen av sista meningen i artikel 12.4 a i konventionen rör i huvudsak två frågor. Den första är huruvida denna bestämmelse innehåller någon skyldighet för de medlemsstater som är parter till konventionen och den andra är vilken räckvidd termerna ”rättigheter ifråga om befordring som garanteras” enligt nationella regler ska anses ha.
När det gäller den första frågan erinrar domstolen inledningsvis om att det i artikel 12.4 a i konventionen föreskrivs att styrelsen, i administrativa frågor, varje år på förslag av skolinspektörsnämnderna ska besluta om behovet av lärarpersonal genom inrättande eller indragning av tjänster. Den ska säkerställa en rättvis fördelning av tjänster mellan medlemsstaterna. Den ska tillsammans med regeringarna lösa frågor angående utnämning eller utstationering av lärare på de olika nivåerna och studievägledare i skolan. Personalen ska behålla de rättigheter i fråga om befordring och pension som garanteras enligt nationella regler.
Det framgår således av nämnda bestämmelses lydelse att – medan de tre första meningarna i bestämmelsen tilldelar styrelsen befogenheter som vid behov ska utövas i samarbete med regeringarna – den tredje meningen är formulerad på ett neutralt sätt genom att fastställa att lärarna har rätt att behålla de rättigheter i fråga om befordring och pension som garanteras enligt nationella regler, utan att specificera vem som ska garantera att lärarna behåller dessa rättigheter.
Det är emellertid uppenbart att nämnda rättigheter inte skulle kunna behållas om de medlemsstater som är parter till konventionen var fria att utforma sina nationella regler och de bestämmelser som reglerar utnämning eller utstationering av sina lärare vid en Europaskola på ett sätt som skulle frånta dessa lärare deras rättigheter under den tid som utnämningen eller utstationeringen avser.
I detta avseende påpekar domstolen att de vid Europaskolorna utnämnda eller utstationerade lärarnas rättigheter i fråga om befordring och pension helt och hållet bestäms av respektive nationella regler och att det följaktligen är omöjligt för styrelsen att garantera att dessa rättigheter behålls när dessa regler inte möjliggör att rättigheterna behålls. Styrelsen är visserligen skyldig att iaktta de nationella reglerna, men det är ändå så att tillämpningen av dessa regler på utnämnda eller utstationerade lärare inte kräver något agerande från styrelsens sida och att det är svårt att tänka sig att styrelsen, med beaktande av att styrelsens befogenheter är begränsade och strikt avgränsade av konventionen, kan åsidosätta lärarnas rättigheter i fråga om befordring och pension enligt nationella regler.
Domstolen konstaterar att under sådana omständigheter skulle Förenade kungarikets tolkning av sista meningen i artikel 12.4 a i konventionen – som innebär att bestämmelsen riktar sig uteslutande till styrelsen i syfte att ålägga den att iaktta de nationella reglerna avseende befordring och pension – frånta bestämmelsen all ändamålsenlig verkan.
I motsats till vad Förenade kungariket har gjort gällande ska denna bestämmelse således tolkas på så sätt att den också för de medlemsstater som är parter till konventionen innebär en skyldighet att garantera att lärarna, under den tid utnämningen eller utstationeringen vid Europaskolorna varar, behåller de rättigheter i fråga om befordring och pension som garanteras enligt nationella regler.
Detta konstaterande motsägs varken av det faktum att artikel 12 i konventionen hör till avdelning II med rubriken ”Skolornas organ”, i vilken anges vilka uppgifter styrelsen ska ha i administrativa frågor, eller av den hänvisning som i artikel 3.2 i konventionen görs till artikel 12 i konventionen.
Även om det står klart att artikel 12 i huvudsak anger vad som åligger styrelsen bör det påpekas att denna artikel, i näst sista meningen i punkt 4 a, också avser ”regeringarna” och att sista meningen i denna bestämmelse, som konstaterats ovan i punkt 42 i denna dom, inte är formulerad på ett sådant sätt att den innebär ett åläggande för styrelsen, utan i stället på ett sådant sätt att den anger en ovillkorlig rättighet för de lärare som är utnämnda eller utstationerade vid Europaskolorna.
Placeringen av denna sista mening förklaras av historiska skäl och av det inneboende samband som finns mellan syftet med denna mening och syftet med den föregående meningen. I stadgan för Europaskolan, som avses i punkt 2 i denna dom, i dess lydelse av den 12 april 1957, var dessa meningar förenade och artikel 12.3 i stadgan föreskrev att styrelsen ”tillsammans med regeringarna [skulle avgöra] frågor om utnämning och utstationering av lärare och skolvärdar på ett sådant sätt att dessa behåller sina rättigheter i fråga om befordring och pension som garanteras enligt nationella regler och får del av de förmåner som tilldelas tjänstemännen i deras kategori i utlandet”. Det framgår tydligt av denna tidigare lydelse av stadgan att styrelsen och regeringarna tillsammans skulle avgöra frågor om utnämning och utstationering på ett sådant sätt att lärarna inte missgynnades på grund av deras utnämning eller utstationering vid en Europaskola. Även om konventionen i sin nuvarande lydelse ytterligare stärker skyddet för lärarna genom att tillerkänna dem en uttrycklig och ovillkorlig rättighet, avser den på intet sätt att befria regeringarna från deras skyldigheter i detta avseende.
I motsats till vad Förenade kungariket tycks anse, är dessutom denna skyldighet inte utan innehåll på grund av det faktum att medlemsstaterna är skyldiga att följa sin egen lagstiftning. Det framgår nämligen ovan att det ansvar som de medlemsstater som är parter till konventionen har för att uppnå det mål som avses i sista meningen i artikel 12.4 a i konventionen inte bara innefattar skyldigheten att iaktta nationella regler i fråga om befordring och pension, utan också skyldigheten att garantera att dessa regler utformas på ett sådant sätt att de inte utesluter lärare som är utnämnda eller utstationerade vid Europaskolorna.
En sådan skyldighet är dessutom inte oförenlig med artikel 165 FEUF. För det första berör den begränsning av Europeiska unionens befogenhet på utbildningsområdet som föreskrivs i denna artikel inte konventionen, eftersom denna inte är en sekundärrättsakt som antagits av ett av unionens organ, utan ett folkrättsligt avtal som ingåtts mellan medlemsstaterna och Europeiska gemenskaperna. Vad för det andra gäller det som anges i tredje skälet i konventionen – att det samarbetssystem av sitt eget slag mellan medlemsstaterna och Europeiska gemenskaperna som det är fråga om erkänner medlemsstaternas ansvar för organisationen av sina utbildningssystem – kan det konstateras att detta ansvar inte på något sätt påverkas av medlemsstaternas skyldighet att inte missgynna de lärare som är utnämnda eller utstationerade vid Europaskolorna i fråga om rättigheter till befordring och pension.
När det gäller den andra tolkningsfrågan – som parterna har olika uppfattning om och som avser vilken räckvidd termerna ”rättigheter ifråga om befordring som garanteras” enligt nationella regler, som återfinns i sista meningen i artikel 12.4 a i konventionen, ska anses ha – bör det påpekas att räckvidden av denna bestämmelse och därigenom det skydd som denna bestämmelse ger de lärare som är utnämnda eller utstationerade vid Europaskolorna inte kan skilja sig åt beroende på varifrån lärarna kommer och att nämnda termer således ska ges en självständig tolkning.
En sådan tolkning måste bland annat göra det möjligt att faktiskt uppnå målet med denna bestämmelse och måste således garantera att lärarna inte missgynnas i fråga om rättigheter till befordring och pension på grund av deras utnämning eller utstationering vid Europaskolorna.
När det gäller termen ”befordring” kan domstolen, mot bakgrund av nämnda mål med bestämmelsen, inte godta den restriktiva tolkning som Förenade kungariket har föreslagit. Såsom generaladvokaten har påpekat i punkterna 45 och 46 i sitt förslag till avgörande, avser denna term inte bara en lärares befordran till tjänster med en högre ställning i en skolas hierarki och som är förknippade med ett större ansvar, såsom en rektorstjänst, utan allt avancemang i karriären. Termen omfattar således även uppflyttning till högre tjänstegrader inom samma befattning, varvid den berörde får högre lön men inte vare sig en annan tjänstebeteckning eller utökat ansvar.
I motsats till vad Förenade kungariket tycks anse går det inte av termerna ”rättigheter som garanteras” enligt nationella regler att sluta sig till att det enda som avses i princip är fall där det i nationella regler föreskrivs en automatisk befordran med koppling till tjänstgöringstid. Såsom generaladvokaten har angett i punkterna 53–55 i sitt förslag till avgörande, framgår det av lydelsen av och ändamålet med den sista meningen i artikel 12.4 a i konventionen att denna bestämmelse avser att se till att lärare som är utnämnda eller utstationerade vid Europaskolorna får behålla alla rättigheter i fråga om karriärutveckling som föreskrivs i respektive nationella regler, oberoende av den form som dessa rättigheter har. Beroende på innehållet i de rättigheter som erkänns i dessa regler kan dessa rättigheter exempelvis innebära en automatisk rätt till befordran eller enbart en rätt att delta i de förfaranden som gör det möjligt att komma vidare i karriären. Däremot kan dessa rättigheter inte vara mer begränsade än de rättigheter som dessa lärare skulle ha åtnjutit om de hade stannat kvar på sin tjänst vid skolan i sin ursprungsmedlemsstat.
Av det ovan anförda följer att artikel 12.4 a sista meningen i konventionen ska tolkas så, att den förpliktar de medlemsstater som är parter till denna konvention att se till att de lärare som är utstationerade eller utnämnda vid Europaskolorna – under den tid som utstationeringen eller utnämningen varar – åtnjuter samma rättigheter i fråga om karriärutveckling och pension som dem som är tillämpliga på deras nationella motsvarigheter enligt deras ursprungsmedlemsstats regler.
Förenade kungarikets tillämpning av artikel 12.4 a sista meningen och artikel 25.1 i konventionen
Parternas argument
Kommissionen anser att det anställningsavtal som engelska och walesiska lärare måste ingå med utbildningsministeriet för deras utstationering vid Europaskolorna är oförenligt med artiklarna 12.4 a och 25.1 i konventionen, eftersom det innebär att lönen för dessa lärare fryses vid då gällande löneklass för hela utstationeringsperioden och eftersom det hindrar dem från att ansöka om att flyttas upp till en högre löneklass eller komma i åtnjutande av de ”teaching and learning responsibility payments” som föreskrivs i STPCD.
Enligt kommissionen missgynnas de potentiella sökandena genom att det är omöjligt för dem att, under den tid utstationeringen varar, delta i den utvärdering som möjliggör för dem att få tillträde till ”post-threshold pay scale”. På grund av detta kan de, när de återvänder till Förenade kungariket efter utstationeringen, endast söka tjänster som omfattas av grundlöneskalan, vilket begränsar utbudet av tillgängliga tjänster.
Det faktum att lärarna i fråga under en nioårig utstationering inte kan komma i fråga för tilläggsbetalningar eller befordringar minskar enligt kommissionen i betydande utsträckning den lön som beaktas vid beräkningen av pensionsrättigheter och således storleken på den framtida pensionen för dessa lärare.
Kommissionen har dessutom gjort gällande att detta har en betydande negativ inverkan på unionens budget, eftersom unionens budget måste täcka en större skillnad mellan den lägre nationella lönen och den harmoniserade lönen enligt stadgan för den utstationerade personalen.
Kommissionen anser, med utgångspunkt i en ungefärlig uträkning, att unionens budget år 2008 var tvungen att täcka extra kostnader på ungefär 720000 euro för de 194 engelska och walesiska utstationerade lärarna. Denna kostnad är resultatet av den större skillnad som måste täckas enligt artikel 49.2 b i stadgan för den utstationerade personalen och följaktligen enligt artikel 25.2 i konventionen. Med utgångspunkt i denna uträkning kan det skäligen anses att det faktum att det är omöjligt för de engelska och walesiska utstationerade lärarna att få tillträde till ”post-threshold pay scale” orsakar en extra årlig kostnad för unionens budget på mellan 500000 och 1000000 euro.
Kommissionen har påpekat att den inte anser att de engelska och walesiska utstationerade lärarna automatiskt måste få tillträde till de högre löneskalorna för ”post-threshold teacher”, ”advanced teacher” och ”excellent teacher” och avancera inom dessa på samma sätt eller få del av ”teaching and learning responsibility payments”. Kommissionen anser det vara tillräckligt att dessa lärare får del av löneutvecklingen på samma villkor som alla andra lärare som är anställda i Förenade kungariket och att de således bland annat kan delta i de utvärderingsförfaranden som föreskrivs för tillträde till dessa löneskalor.
Enligt kommissionen framgår det av en noggrann undersökning av de olika yrkesmässiga normer och uppgifter som gäller avseende dessa löneskalor och tilläggsbetalningar att de lärare som är utstationerade vid Europaskolorna utför sådana uppgifter som i princip är ägnade att ge dem tillträde till nämnda löneskalor eller få del av nämnda tilläggsbetalningar.
Kommissionen anser att Förenade kungariket inte kan åberopa påstådda tekniska svårigheter för att rättfärdiga åsidosättandet av de skyldigheter som följer av konventionen. Dessutom ifrågasätter kommissionen att sådana svårigheter faktiskt föreligger eller att dessa svårigheter inte skulle kunna överbryggas med hjälp av insatser som står i proportion till de intressen som berörs.
När det för det första gäller genomförandet av utvärderingen av de utstationerade lärarna, har kommissionen påpekat att utvärderingen avseende tillträde till ”post-threshold pay scale” utförs av rektorerna vid respektive skola och att det inte tycks finnas något som hindrar att denna uppgift anförtros rektorn vid Europaskolan. Även andra lösningar är tänkbara. Förenade kungariket skulle kunna sända inspektörer som kontrollerar den utvärdering som rektorerna vid Europaskolorna genomför. Utvärderingen skulle kunna genomföras av utomstående. Även en kombination av dessa båda lösningar är tänkbar. Slutligen finns det inget som hindrar att de utvärderare från den nationella myndigheten som utför utvärderingarna av nationella sökande till ”advanced skills teachers”- och ”excellent teachers”-tjänsterna kommer till Europaskolorna, eftersom de redan utför utvärderingar i försvarsministeriets skolor i Tyskland och i andra länder utanför Förenade kungariket.
När det för det andra gäller Förenade kungarikets argument som grundar sig på att tillträdet till högre löneskalor är beroende av inrättandet av tjänster, har kommissionen påpekat att detta inte är fallet när det gäller tillträde till ”post-threshold pay scale”, vars införande i huvudsak utgör en förtäckt generell lönehöjning. När det gäller tillträdet till övriga högre löneskalor rör det sig om att skapa en tjänst i budgethänseende. Emellertid finns det inget som hindrar Förenade kungariket från att tilldela utbildningsministeriet ett lämpligt antal ”advanced skills teachers”- och ”excellent teachers”-tjänster för de utstationerade lärarna.
Förenade kungariket har ifrågasatt påståendet att dess behandling av de utstationerade lärarna strider mot artiklarna 12.4 a och 25 i konventionen.
Förenade kungariket anser att kommissionens talan bygger på en felaktig förståelse av stadgan för de utstationerade lärarna och av karaktären av de tilläggsbetalningar som föreskrivs i STPCD. I detta avseende har denna medlemsstat bland annat påpekat att de engelska och walesiska utstationerade lärarna inte nödvändigtvis tidigare var verksamma vid en nationell statsunderstödd skola och därför inte nödvändigtvis omfattades av STPCD före utstationeringen. STPCD utgör därför inte de ”nationella regler[na]” i den mening som avses i artikel 12 i konventionen.
Enligt Förenade kungariket har dessutom de utstationerade engelska och walesiska lärarna frivilligt lämnat sina tidigare tjänster för en ny tjänst vid en Europaskola på grundval av ett nytt anställningskontrakt som ingåtts med utbildningsministeriet. I nämnda kontrakt anges också att en utstationerad lärare inte kan ansöka om att få tillträde till de högre löneskalorna och de tilläggsbetalningar som avses i STPCD. Nämnda lärare har således frivilligt valt en tjänst som inte omfattas av STPCD.
För övrigt har Förenade kungariket gjort gällande att de tilläggsbetalningar som föreskrivs i STPCD inte ”garanteras” enligt nationella regler och inte utgör ”rättigheter i fråga om befordring”, i den mening som avses i artikel 12.4 a i konventionen. Dessa tilläggsbetalningar följer inte automatiskt av tjänstgöringstid, utan läraren måste ansöka om dem, och de tilldelas endast enligt vissa villkor. Dessutom är ”teaching and learning responsibility payments” och ”advanced skills teachers”- och ”excellent teachers”-systemen endast tillgängliga för det fall en skola beslutar att inrätta sådana tjänster. Tilläggsbetalningarna utgör inte heller en ”befordring” i den mening som avses i nämnda artikel, eftersom de lärare som får en sådan betalning fortfarande tjänstgör som ”lärare” och inte får en högre uppsatt tjänst.
Förenade kungariket anser att om de utstationerade lärarna hade rätt till tilläggsbetalningar utan att behöva utöva det ansvar som är förknippat med dem, skulle detta innebära att de lärare som är verksamma i Förenade kungariket diskriminerades. Förenade kungariket har bland annat bestritt att de utstationerade lärarna uppfyller de villkor som uppställs för att de ska få tilläggsbetalningar. Således föreligger inte någon faktisk likvärdighet mellan situationen för de europeiska lärarna och situationen för lärarna vid de statsunderstödda skolorna i Förenade kungariket.
Enligt Förenade kungariket skulle det faktum att kontrollen av Europaskolornas lärares yrkesmässiga kompetens inte skulle vara lika noggrann och sträng som den kontroll som föreskrivs på nationell nivå även utgöra en diskriminering av de lärare som är verksamma i Förenade kungariket. Den lösning som kommissionen föreslår – att nämnda kontroll utförs av inspektörer som utsänds från Förenade kungariket vid Europaskolorna – är inte tillräcklig för att garantera en likvärdighet i detta avseende.
När det slutligen gäller artikel 25 i konventionen har Förenade kungariket gjort gällande att även om Förenade kungarikets tolkning av artikel 12.4 a sista meningen i konventionen visade sig vara felaktig, skulle det ändå inte föreligga någon förlust för unionens budget. Det är visserligen möjligt att en del av de utstationerade och utnämnda engelska och walesiska lärarna vid Europaskolorna förvärvar rätten att få del av en tilläggsbetalning i framtiden, om de ger in en lämplig ansökan och denna godkänns. Eftersom beviljandet av en sådan rättighet är beroende av en individuell utvärdering av varje lärare, kan emellertid för närvarande inte någon av nämnda lärare göra anspråk på en sådan. Följaktligen har Förenade kungariket hittills fullgjort sin skyldighet att betala hela beloppet avseende lön som dessa lärare har rätt till.
Domstolens bedömning
Kommissionen har i huvudsak gjort gällande att Förenade kungariket har underlåtit att i enlighet med artikel 12.4 a sista meningen i konventionen se till att de lärare som England och Wales har utnämnt eller utstationerat vid Europaskolorna får behålla de rättigheter i fråga om befordring och pension som garanteras enligt nationella regler och följaktligen också, i strid med artikel 25.1 i samma konvention, underlåtit att fortsätta att betala ut lön till dessa lärare.
För att bedöma huruvida detta påstående är välgrundat prövar domstolen först huruvida STPCD för dessa lärare utgör de nationella regler som gäller för lärarna i fråga, i den mening som avses i artikel 12.4 a sista meningen i konventionen.
I detta avseende är det av betydelse att pröva huruvida medlemsstaterna som är parter till konventionen – även om de, såsom det erinras om i tredje skälet i konventionen, fortfarande är helt och hållet ansvariga för organisationen av sina utbildningssystem – är förhindrade att åberopa särdrag i utbildningssystemet för att undandra sig skyldigheter som följer av konventionen och för att frånta de lärare som de utnämner eller utstationerar vid Europaskolorna det skydd som föreskrivs i artikel 12.4 a sista meningen i konventionen.
Detta skulle vara följden av Förenade kungarikets argumentation som går ut på att STPCD inte utgör de nationella reglerna för de engelska och walesiska lärarna i den mening som avses i nämnda bestämmelse. Enligt denna argumentation skulle det, med beaktande av särdragen i denna medlemsstats utbildningssystem, helt enkelt inte finnas några nationella regler för den medlemsstaten.
Dessutom bör det påpekas att STPCD är obligatoriskt för alla statsunderstödda skolor i England och Wales och att majoriteten av de lärare som anställs inom dessa områden är anställda av en sådan skola. Påpekas bör även den omständigheten att också en stor del av de icke-statsunderstödda skolorna helt eller delvis tillämpar STPCD. Kommissionen har i detta avseende anfört, utan att på denna punkt bli motsagd av Förenade kungariket, att de icke-statsunderstödda skolor som endast delvis tillämpar STPCD i praktiken använder sig av de villkor som föreskrivs i STPCD som utgångspunkt och lägger till ytterligare förmåner samt att STPCD i själva verket tillämpas på 90 procent av de lärare som är anställda i denna medlemsstat.
Det standardanställningsavtal, som de lärare som är utnämnda eller utstationerade av England och Wales vid Europaskolorna ingår med utbildningsministeriet med anledning av utnämningen eller utstationeringen, föreskriver dessutom att de nationella löner som varje månad betalas ut till dessa lärare ska fastställas i enlighet med löneskalorna i STPCD och att dessa lärare ska ha rätt till årliga löneökningar som förhandlas fram på nationell nivå och är tillämpliga i kraft av STPCD. Det står således klart att även för nämnda lärare är arbetsförhållandena delvis reglerade genom STPCD och att det alltså endast är selektivt, bland annat när det gäller möjligheten till en högre löneskala och en tilläggsbetalning, som nämnda avtal utesluter tillämpningen av STPCD.
Vid dessa förhållanden måste det konstateras att STPCD utgör de nationella reglerna för de engelska och walesiska lärarna i den mening som avses i artikel 12.4 a sista meningen i konventionen.
När det gäller Förenade kungarikets argument att Förenade kungariket inte är skyldigt att tillerkänna alla de lärare som det utnämner eller utstationerar vid Europaskolorna de rättigheter i fråga om befordring som föreskrivs i STPCD, eftersom endast en del av dessa lärare före utnämningen eller utstationeringen var verksamma vid en statsunderstödd skola i England eller Wales, bör det påpekas att kommissionen inom ramen för denna talan inte har påstått att nämnda i STPCD föreskrivna rättigheter ska tillämpas på alla lärare som Förenade kungariket har utnämnt eller utstationerat, utan endast på de lärare som kommer från England och Wales. Den omständigheten att STPCD bland annat inte tillämpas på de lärare som är anställda i Skottland saknar följaktligen betydelse för prövningen av denna talan.
I den mån som inte bara de statsunderstödda skolorna i England och Wales, utan också en stor andel av de icke-statsunderstödda skolorna, helt eller delvis tillämpar STPCD, kan det för övrigt antas att flertalet av de engelska och walesiska utnämnda eller utstationerade lärarna vid Europaskolorna omfattades av villkoren i STPCD före utnämningen eller utstationeringen. Även om det skulle visa sig att en del av dessa lärare inte omfattades av STPCD på grund av att de antingen var anställda vid en icke-statsunderstödd skola som inte frivilligt tillämpade STPCD eller inte anställda vid någon skola alls, kan denna omständighet i vilket fall som helst inte motivera att Förenade kungariket, med stöd av det standardavtal som lärarna måste ingå med anledning av utnämningen eller utstationeringen vid Europaskolorna, utesluter samtliga engelska och walesiska lärare från vissa förmåner som föreskrivs i STPCD.
I motsats till vad Förenade kungariket har gjort gällande, motiveras denna uteslutning inte av det faktum att nämnda lärare undertecknar detta avtal med fri vilja och full insikt. Förvisso är det så att dessa lärare inte på något sätt är tvungna att ansöka om att utnämnas eller utstationeras vid en Europaskola samt kan ta reda på innehållet i det nya anställningsavtalet. Dessa lärare har dock inget annat val än att underteckna nämnda avtal, vars villkor påtvingas dem av utbildningsministeriet. Utan att frånta artikel 12.4 a sista meningen i konventionen dess ändamålsenliga verkan kan det under sådana omständigheter inte på goda grunder anses att lärarna frivilligt har avstått från nämnda i STPCD föreskrivna förmåner och de rättigheter som de tillerkänns i denna bestämmelse i konventionen.
Domstolen prövar därefter frågan huruvida tillträdet till mer fördelaktiga löneskalor, såsom ”post-threshold pay scale” och de löneskalor som tillämpas på ”excellent teachers” och ”advanced skills teachers”, samt åtnjutandet av andra tilläggsbetalningar, såsom ”teaching and learning responsibility payments”, som föreskrivs i STPCD, utgör rättigheter i fråga om befordring, i den mening som avses i den bestämmelsen. I detta avseende erinrar domstolen om att det redan har konstaterats i punkterna 54 och 55 i denna dom att även sådana rättigheter som innebär högre lön men inte en annan tjänstebeteckning för läraren, liksom sådana rättigheter som inte automatiskt tilldelas på grundval av tjänstgöringstid utan kräver att läraren deltar i förfaranden och uppfyller vissa villkor, utgör rättigheter i fråga om befordring, i den mening som avses i den bestämmelsen.
Av detta följer att domstolen inte kan godta Förenade kungarikets argument att de lärare, för vilka dessa löneskalor och betalningar gäller, har behållit sina befattningar och har behövt underkasta sig sådana förfaranden. Dessutom har kommissionen inte gjort gällande att de lärare som är utnämnda eller utstationerade av England eller Wales automatiskt måste få del av nämnda löneskalor och betalningar, men att de måste ha tillgång till dem på samma villkor som dem som gäller för engelska och walesiska lärare som omfattas av STPCD.
Förenade kungariket har gjort gällande att de utnämnda eller utstationerade lärarna i princip inte kan uppfylla de yrkesmässiga normer som måste vara uppfyllda för att en lärare ska få tillträde till dessa löneskalor samt utöva sådant ytterligare ansvar som är kopplat till tillämpningen av vissa av dessa löneskalor och betalningar. Domstolen påpekar i detta avseende att kommissionen har gjort en noggrann undersökning av dessa krav och åtaganden och därvid på ett rimligt sätt förklarat att ett stort antal av nämnda lärare uppfyller dessa normer och har likvärdiga åtaganden vid Europaskolorna.
Denna undersökning och dessa förklaringar har inte ifrågasatts genom de enstaka argument som framförts av Förenade kungariket och som i huvudsak går ut på att det inte föreligger någon faktisk likvärdighet mellan situationen för lärarna vid Europaskolorna och situationen för deras nationella motsvarigheter. Ett sådant påstående strider faktiskt mot artikel 10 i stadgan för den utstationerade personalen, enligt vilken de utnämnda eller utstationerade lärarna ska besitta de kvalifikationer och uppfylla de nödvändiga villkor som erfordras för att inneha motsvarande befattningar i de länder de kommer från. I den mån som nämnda argument grundar sig på uppfattningen att nämnda lärare per definition inte kan uppfylla dessa normer och ha sådana åtaganden mot bakgrund av att Europaskolorna inte fungerar exakt likadant som de statsunderstödda skolorna i England och Wales, beaktar inte argumenten Europaskolornas särskilda ställning och att de utgör ett system av sitt eget slag.
I motsats till vad Förenade kungariket har gjort gällande, innebär tillträdet till nämnda löneskalor och tilläggsbetalningar för de lärare som är utnämnda eller utstationerade av England och Wales vid Europaskolorna inte heller en diskriminering av deras nationella motsvarigheter med hänvisning till att det är omöjligt att utföra kontroller av Europaskolornas lärares yrkesmässiga kompetens lika noggrant och strängt som kontrollerna på nationell nivå. Såsom generaladvokaten har påpekat i punkterna 87–90 i sitt förslag till avgörande, är detta argument ogrundat, eftersom det är helt och hållet genomförbart att utföra sådana kontroller. Förenade kungariket har för övrigt inte närmare angett varför det anser att de olika lösningar som i detta avseende har föreslagets av kommissionen inte möjliggör att ett tillfredsställande resultat uppnås, utan har inskränkt sig till att påstå att det inte skulle vara tillräckligt att skicka nationella inspektörer till Europaskolorna.
Förenade kungariket har också anfört att många lärare vid de statsunderstödda skolorna i England och Wales inte omfattas av de löneskalor som föreskrivs för ”excellent teachers” och ”advanced skills teachers” eller ”teaching and learning responsibility payments” på grund av att ingen sådan tjänst eller mycket få sådana tjänster som ger rätt till dessa löneskalor och betalningar har inrättats vid deras skolor. Denna omständighet motiverar emellertid inte att samtliga engelska och walesiska utnämnda eller utstationerade lärare vid Europaskolorna utesluts från dessa löneskalor och betalningar.
Som svar på kommissionens begäran om inrättande vid Europaskolorna av ett antal sådana tjänster som står i proportion till antalet i England och Wales, har Förenade kungariket inte ifrågasatt att detta faktiskt är möjligt, men har uppgett att det antal tjänster som skulle inrättas vid Europaskolorna skulle vara mycket lågt eller till och med obefintligt och att det vid dessa förhållanden skulle vara svårt att avgöra vid vilka Europaskolor dessa tjänster skulle inrättas. Sådana praktiska svårigheter vid fördelningen av tjänster som ger rätt till nämnda löneskalor och betalningar kan emellertid inte motivera att några sådana tjänster inte inrättas vid Europaskolorna. Det står dessutom klart att Förenade kungariket, med stöd av artikel 12.4 a näst sista meningen i konventionen, kan få hjälp av styrelsen med att lösa dessa problem för att bland annat identifiera tjänster vid Europaskolorna att besätta med ”excellent teachers” och ”advanced skills teachers”.
Av det ovan anförda framgår att tillträdet till mer fördelaktiga löneskalor, såsom ”post-threshold pay scale” och de löneskalor som tillämpas på ”excellent teachers” och ”advanced skills teachers”, samt åtnjutandet av andra tilläggsbetalningar, såsom ”teaching and learning responsibility payments”, som föreskrivs i STPCD, utgör rättigheter i fråga om befordring, i den mening som avses i artikel 12.4 a sista meningen i konventionen, vilka Förenade kungariket måste säkerställa att de lärare som England och Wales har utnämnt eller utstationerat vid Europaskolorna omfattas av. Eftersom tillträdet till dessa löneskalor och betalningar har en direkt påverkan på storleken på den pension som dessa lärare kan kräva, utgör dessa också en rättighet i fråga om pension som garanteras enligt nationella regler i den mening som avses i den bestämmelsen.
När det slutligen gäller frågan huruvida Förenade kungariket tillämpar artikel 25.1 i konventionen korrekt, erinrar domstolen om att denna bestämmelse ålägger medlemsstaterna att bidra till Europaskolornas budget genom bidrag i form av fortsatt utbetalning av lön till de lärare som de utstationerar eller utnämner vid dessa skolor. Enligt punkt 2 i samma artikel, jämförd med artikel 49 i stadgan för den utstationerade personalen, ska unionen bidra till nämnda budget genom att betala det europeiska tillägget. I detta avseende har kommissionen, utan att bli motsagd av Förenade kungariket på denna punkt, företett sifferuppgifter som på ett rimligt sätt visar att frysningen av lönerna för de engelska och walesiska lärare som är utnämnda eller utstationerade vid Europaskolorna har gjort att unionen har varit tvungen att betala ett högre europeiskt tillägg till dessa lärare, vilket har orsakat en ökning av unionens årliga bidrag till skolornas budget.
Denna bedömning påverkas inte av Förenade kungarikets argument att tillträdet till de högre löneskalorna och tilläggsbetalningarna är beroende av en individuell utvärdering av varje lärare, vilken fortfarande inte har gjorts avseende de engelska och walesiska lärare som är utnämnda eller utstationerade vid Europaskolorna. Detta argument beaktar uppenbarligen inte vare sig att anledningen till att dessa utvärderingar inte ägt rum är att dessa lärare systematiskt har uteslutits från nämnda löneskalor och betalningar eller det faktum att det rimligen kan antas att vissa av dessa lärare redan skulle ha fått tillträde till dessa löneskalor och betalningar om de inte varit uteslutna därifrån.
Av detta följer att i den mån som en korrekt tolkning och en korrekt tillämpning av Förenade kungariket av artikel 12.4 a sista meningen i konventionen skulle ha lett till att denna medlemsstat bidrog i större utsträckning till Europaskolornas budget, finns det ett åtminstone indirekt samband mellan åsidosättandet av artikel 12.4 a i konventionen och den skyldighet som åligger medlemsstaterna enligt artikel 25.1 i konventionen. Detta samband har för övrigt inte bestritts av Förenade kungariket. Följaktligen har Förenade kungariket, genom att hindra nämnda lärare från att ansöka om att omfattas av en högre löneklass eller komma i åtnjutande av ”teaching and learning responsibility payments”, också åsidosatt artikel 25.1 i konventionen.
Mot bakgrund av det ovan anförda konstaterar domstolen följande. Förenade kungariket har gjort en felaktig tillämpning av artiklarna 12.4 a och 25.1 i konventionen genom att utesluta de engelska och walesiska lärare som är utnämnda eller utstationerade vid Europaskolorna, under den tid som utnämningen eller utstationeringen varar, från tillträde till mer fördelaktiga löneskalor, bland annat ”threshold pay”, ”excellent teacher system” och ”advanced skills teachers” och tillträde till andra i STPCD föreskrivna tilläggsbetalningar, såsom ”teaching and learning responsibility payments”.
Rättegångskostnader
Enligt artikel 69.2 i rättegångsreglerna ska tappande part förpliktas att ersätta rättegångskostnaderna, om detta har yrkats. Kommissionen har yrkat att Förenade kungariket ska förpliktas att ersätta rättegångskostnaderna. Eftersom Förenade kungariket har tappat målet, ska kommissionens yrkande bifallas.
Mot denna bakgrund beslutar
domstolen (första avdelningen)
följande:
Artikel 12.4 a sista meningen i konventionen med stadga för Europaskolorna av den 21 juni 1994 ska tolkas så, att den förpliktar de medlemsstater som är parter till denna konvention att se till att de lärare som är utstationerade eller utnämnda vid Europaskolorna – under den tid som utstationeringen eller utnämningen varar – åtnjuter samma rättigheter i fråga om karriärutveckling och pension som dem som är tillämpliga på deras nationella motsvarigheter enligt deras ursprungsmedlemsstats regler.
Förenade konungariket Storbritannien och Nordirland har gjort en felaktig tillämpning av artiklarna 12.4 a och 25.1 i konventionen genom att utesluta de engelska och walesiska lärare som är utnämnda eller utstationerade vid Europaskolorna, under den tid som utnämningen eller utstationeringen varar, från tillträde till mer fördelaktiga löneskalor, bland annat ”threshold pay”, ”excellent teacher system” och ”advanced skills teachers” och tillträde till andra i ”School Teachers Pay and Conditions Document” föreskrivna tilläggsbetalningar, såsom ”teaching and learning responsibility payments”.
Förenade konungariket Storbritannien och Nordirland ska ersätta rättegångskostnaderna.
Underskrifter
Artikel 267 FEUF — Upphävande av ett domstolsavgörande — Återförvisning till berörd domstol — Skyldighet att följa beslutet om upphävande — Begäran om förhandsavgörande — Möjlighet — Miljö — Århuskonventionen — Direktiv 85/337/EEG — Direktiv 96/61/EG — Allmänhetens deltagande i beslutsprocesser — Anläggande av en avfallsdeponi — Ansökan om tillstånd — Affärshemligheter — En handling har inte gjorts tillgänglig för allmänheten — Verkningar för giltigheten av beslutet att meddela tillstånd för deponin — Rättelse — Miljökonsekvensbedömning av projektet — Slutligt utlåtande har utfärdats före medlemsstatens anslutning till unionen — Tillämplighet i tiden av direktiv 85/337 — Rättsmedel — Interimistiska åtgärder — Inhibition — Upphävande av det angripna beslutet — Äganderätt — Ingrepp”
I mål C-416/10,
angående en begäran om förhandsavgörande enligt artikel 267 FEUF, framställd av Najvyšší súd Slovenskej republiky (Slovakien) genom beslut av den 17 augusti 2010, som inkom till domstolen den 23 augusti 2010, i målet
Jozef Križan,
Katarína Aksamitová,
Gabriela Kokošková,
Jozef Kokoška,
Martina Strezenická,
Jozef Strezenický,
Peter Šidlo,
Lenka Šidlová,
Drahoslava Šidlová,
Milan Šimovič,
Elena Šimovičová,
Stanislav Aksamit,
Tomáš Pitoňák,
Petra Pitoňáková,
Mária Križanová,
Vladimír Mizerák,
Ľubomír Pevný,
Darina Brunovská,
Mária Fišerová,
Lenka Fišerová,
Peter Zvolenský,
Katarína Zvolenská,
Kamila Mizeráková,
Anna Konfráterová,
Milan Konfráter,
Michaela Konfráterová,
Tomáš Pavlovič,
Jozef Krivošík,
Ema Krivošíková,
Eva Pavlovičová,
Jaroslav Pavlovič,
Pavol Šipoš,
Martina Šipošová,
Jozefína Šipošová,
Zuzana Šipošová,
Ivan Čaputa,
Zuzana Čaputová,
Štefan Strapák,
Katarína Strapáková,
František Slezák,
Agnesa Slezáková,
Vincent Zimka,
Elena Zimková,
Marián Šipoš,
Mesto Pezinok
mot
Slovenská inšpekcia životného prostredia,
ytterligare deltagare i rättegången:
Ekologická skládka as,
meddelar
DOMSTOLEN (stora avdelningen)
sammansatt av ordföranden V. Skouris, vice ordföranden K. Lenaerts, avdelningsordförandena A. Tizzano, M. Ilešič, L. Bay Larsen (referent) och J. Malenovský samt domarna A. Borg Barthet, J.-C. Bonichot, C. Toader, J.-J. Kasel och M. Safjan,
generaladvokat: J. Kokott,
justitiesekreterare: handläggaren C. Strömholm,
efter det skriftliga förfarandet och förhandlingen den 17 januari 2012,
med beaktande av de yttranden som avgetts av:
Jozef Križan, Katarína Aksamitová, Gabriela Kokošková, Jozef Kokoška, Martina Strezenická, Jozef Strezenický, Peter Šidlo, Lenka Šidlová, Drahoslava Šidlová, Milano Šimovič, Elena Šimovičová, Stanislav Aksamit, Tomáš Pitoňák, Petra Pitoňáková, Mária Križanová, Vladimír Mizerák, Ľubomír Pevný, Darina Brunovská, Mária Fišerová, Lenka Fišerová, Peter Zvolenský, Katarína Zvolenská, Kamila Mizeráková, Anna Konfráterová, Milano Konfráter, Michaela Konfráterová, Tomáš Pavlovič, Jozef Krivošík, Ema Krivošíková, Eva Pavlovičová, Jaroslav Pavlovič, Pavol Šipoš, Martina Šipošová, Jozefína Šipošová, Zuzana Šipošová, Ivan Čaputa, Zuzana Čaputová, Štefan Strapák, Katarína Strapáková, František Slezák, Agnesa Slezáková, Vincent Zimka, Elena Zimková och Marián Šipoš, genom T. Kamenec och Z. Čaputová, advokáti,
Mesto Pezinok, genom J. Ondruš och K. Siváková, advokáti,
Slovenská inšpekcia životného prostredia, genom L. Fogaš, advokát,
Ekologická skládka as, genom P. Kováč, advokát,
Slovakiens regering, genom B. Ricziová, i egenskap av ombud,
Tjeckiens regering, genom M. Smolek och. D. Hadroušek, båda i egenskap av ombud,
Frankrikes regering, genom S. Menez, i egenskap av ombud,
Österrikes regering, genom C. Pesendorfer, i egenskap av ombud,
Europeiska kommissionen, genom P. Oliver och A. Tokár, båda i egenskap av ombud,
och efter att den 19 april 2012 ha hört generaladvokatens förslag till avgörande,
följande
Dom
Begäran om förhandsavgörande avser tolkningen av konventionen om tillgång till information, allmänhetens deltagande i beslutsprocesser och tillgång till rättslig prövning i miljöfrågor, som undertecknades i Århus den 25 juni 1998 och som godkändes på Europeiska gemenskapens vägnar genom rådets beslut 2005/370/EG av den 17 februari 2005 (EUT L 124, s. 1) (nedan kallad Århuskonventionen), av artiklarna 191.1 FEUF, 191.2 FEUF och 267 FEUF och av rådets direktiv 85/337/EEG av den 27 juni 1985 om bedömning av inverkan på miljön av vissa offentliga och privata projekt (EGT L 175, s. 40 ; svensk specialutgåva, område 15, volym 6, s. 226), i dess lydelse enligt Europaparlamentets och rådets direktiv 2003/35/EG av den 26 maj 2003 (EUT L 156, s. 17) (nedan kallat direktiv 85/337) samt av rådets direktiv 96/61/EG av den 24 september 1996 om samordnade åtgärder för att förebygga och begränsa föroreningar (EGT L 257, s. 26), i dess lydelse enligt Europaparlamentets och rådets förordning (EG) nr 166/2006 av den 18 januari 2006 (EUT L 33, s. 1) (nedan kallat direktiv 96/61).
Begäran har framställts i ett mål mellan, å ena sidan, Jozef Križan och 43 andra fysiska personer boende i staden Pezinok samt Mesto Pezinok (Pezinok stad) och, å andra sidan, Slovenská inšpekcia životného prostredia (den slovakiska miljöinspektionen) (nedan kallad Inšpekcia) avseende lagenligheten av de myndighetsbeslut varigenom Ekologická skládka as (nedan kallat Ekologická skládka), som intervenerat i det nationella målet, beviljats tillstånd att anlägga och driva en avfallsdeponi.
Tillämpliga bestämmelser
Internationell rätt
I punkterna 1, 2, 4 och 6 i artikel 6 i Århuskonventionen, som har rubriken ”Allmänhetens deltagande i beslut om vissa verksamheter”, föreskrivs följande:
1.   Varje part
skall tillämpa bestämmelserna i denna artikel i fråga om beslut om huruvida sådana föreslagna verksamheter som anges i bilaga I skall tillåtas,
...
I beslutsprocesser om miljön skall den berörda allmänheten på ett tidigt och lämpligt stadium informeras på ett effektivt sätt, antingen genom offentligt tillkännagivande eller i förekommande fall enskilt, bl.a. om:
...
den tänkta beslutsprocessen, inbegripet, om sådan information kan lämnas, information om
...
till vilken myndighet man kan vända sig för att få relevant information och var sådan information finns tillgänglig för allmänhetens granskning,
...
Varje part skall sörja för att allmänhetens deltagande sker på ett tidigt stadium, när alla alternativ är möjliga och allmänheten kan delta på ett meningsfullt sätt.
...
Varje part skall kräva att de behöriga myndigheterna, på begäran när detta krävs enligt nationell rätt, ger den berörda allmänheten möjlighet att kostnadsfritt och så snart informationen blir tillgänglig ta del av all information som är av betydelse för den beslutsprocess som avses i denna artikel och som finns tillgänglig under den tid förfarandet för allmänhetens medverkan pågår, vilket dock inte skall påverka parternas rätt att vägra att lämna ut vissa uppgifter i enlighet med [särskilt artikel 4.4].
...”
I punkterna 2 och 4 i artikel 9 i konventionen, som har rubriken ”Tillgång till rättslig prövning”, föreskrivs följande:
2.   Varje part skall inom ramen för sin nationella lagstiftning se till att den berörda allmänhet[en]
...
... har rätt att få den materiella och formella giltigheten av ett beslut, en handling eller en underlåtenhet som omfattas av artikel 6 eller, om detta föreskrivs i nationell rätt och utan att det påverkar tillämpningen av punkt 3, andra tillämpliga bestämmelser i denna konvention prövad av domstol eller något annat oberoende och opartiskt organ som inrättats genom lag.
...
De förfaranden som avses i punkterna 1–3 skall, utan att det påverkar tillämpningen av punkt 1, erbjuda tillräckliga och effektiva rättsmedel, inbegripet förelägganden där så är lämpligt, och vara objektiva, rättvisa, snabba och inte oöverkomligt kostsamma. …”
I punkt 5 i bilaga I till Århuskonventionen anges, såsom verksamheter som avses i artikel 6.1 a i konventionen, följande:
Avfallshantering:
...
Deponier som tar emot mer än 10 ton avfall per dygn eller med en total kapacitet som överstiger 25000 ton, med undantag för deponier för inert avfall.”
Unionsrätten
Direktiv 85/337
I artikel 1.2 i direktiv 85/337 definieras begreppet ”tillstånd” som ”den ansvariga myndighetens eller de ansvariga myndigheternas beslut, som ger exploatören rätt att genomföra projektet”.
I artikel 2 i direktivet föreskrivs följande:
1.   Medlemsstaterna skall vidta alla nödvändiga åtgärder för att säkerställa att projekt som kan antas medföra en betydande miljöpåverkan bland annat på grund av sin art, storlek eller lokalisering blir föremål för krav på tillstånd och en bedömning av deras påverkan innan tillstånd ges. Dessa projekt anges i artikel 4.
Bedömningen av miljöpåverkan kan integreras i det befintliga tillståndsförfarandet för projekt i medlemsstaterna eller, om detta inte är möjligt, i andra förfaranden eller i sådana förfaranden som tillskapas för att målsättningarna i detta direktiv skall uppfyllas.
...”
Direktiv 96/61
I skäl 23 i direktiv 96/61 föreskrivs följande:
För att allmänhet[en] skall kunna få information om driften vid anläggningarna och dessas eventuella miljöpåverkan och för att säkerställa insynen i tillståndsförfarandena i hela gemenskapen, bör information som rör tillståndsansökningar rörande nya anläggningar… vara tillgängliga för allmänheten [innan något beslut fattas].”
I artikel 1 i direktivet, som har rubriken ”Syfte och tillämpningsområde”, föreskrivs följande:
Detta direktiv syftar till att genom samordnade åtgärder förebygga och minska föroreningar som härrör från de verksamheter som anges i bilaga I. Det innehåller bestämmelser som syftar till att undvika och, när detta visar sig vara omöjligt, minska utsläppen till luft, vatten och mark från dessa verksamheter, inbegripet åtgärder som gäller avfall, så att en hög skyddsnivå kan uppnås för miljön som helhet, utan att detta påverkar tillämpning av bestämmelserna i direktiv [85/337] och andra gemenskapsbestämmelser i ämnet.”
I artikel 15 i direktivet, som har rubriken ”Tillgång till information och allmänhetens deltagande i tillståndsförfarandet”, föreskrivs följande:
1.   Medlemsstaterna skall se till att den berörda allmänheten på ett tidigt stadium ges tillfälle att på ett effektivt sätt deltaga i förfaranden för
meddelande av tillstånd för nya anläggningar,
...
Det förfarande som anges i bilaga V skall tillämpas för sådant deltagande.
...
[Särskilt punkt 1] skall tillämpas med de begränsningar som fastställs i artikel 3.2 och 3.3 i [rådets] direktiv 90/313/EEG [av den 7 juni 1990 om rätt att ta del av miljöinformation (EGT L 158, s. 56; svensk specialutgåva, område 15, volym 9, s. 233)].
...”
I artikel 15a i direktiv 96/61, som har rubriken ”Rätt till rättslig prövning”, föreskrivs följande:
Medlemsstaterna skall inom ramen för den relevanta nationella lagstiftningen se till att … medlemmar[na] av den berörda allmänheten
...
har rätt att få den materiella eller formella giltigheten av ett beslut, en handling eller en underlåtenhet som omfattas av bestämmelserna om allmänhetens deltagande i detta direktiv prövad i domstol eller något annat oberoende och opartiskt organ som inrättats genom lag.
...
Sådana förfaranden skall vara rättvisa, snabba och inte oöverkomligt kostsamma.
...”
I punkt 5.4 i bilaga I till direktiv 96/61, som har rubriken ”Kategorier av industriell verksamhet [som avses i artikel 1]”, hänvisas till ”[a]vfallsdeponier som tar emot mer än 10 ton per dygn eller med en totalkapacitet på mer än 25000 ton, med undantag för avfallsdeponier för inert avfall”.
I bilaga V till direktivet, som har rubriken ”Allmänhetens deltagande i beslutsprocesser”, föreskrivs bland annat följande:
1.
Allmänheten skall informeras (genom offentliga meddelanden eller på annat lämpligt sätt, t.ex. med hjälp av elektroniska medier när sådana är tillgängliga) om följande på ett tidigt stadium under beslutsprocessen och senast så snart som information rimligen kan ges:
...
Uppgifter om vilka myndigheter som är behöriga att fatta beslut, från vilka [myndigheter] relevant information kan erhållas och till [vilka myndigheter] synpunkter eller frågor kan lämnas in samt om tidsfristerna för att överlämna synpunkter eller frågor.
...
Uppgift om när och var eller på vilket sätt relevant information kommer att göras tillgänglig.
...”
Direktiv 2003/4/EG
I skäl 16 i Europaparlamentets och rådets direktiv 2003/4/EG av den 28 januari 2003 om allmänhetens tillgång till miljöinformation och om upphävande av direktiv 90/313 (EUT L 41, s. 26) anges följande:
Rätten till information innebär att den allmänna regeln bör vara att informationen lämnas ut och att offentliga myndigheter bör ha rätt att avslå en begäran om miljöinformation endast i specifika och klart definierade fall. Skälen för avslag bör tolkas restriktivt, varvid allmänhetens intresse av att informationen lämnas ut bör vägas mot det intresse som betjänas av att begäran avslås. Skälen för ett avslag bör vara den sökande tillhanda inom den tidsgräns som fastställs i detta direktiv.”
I artikel 4.2 och 4.4 i direktivet föreskrivs bland annat följande:
2.   Medlemsstaterna får föreskriva att begäran om miljöinformation skall avslås, om utlämnande av informationen skulle ha negativa följder för följande:
...
Sekretess som omfattar kommersiell eller industriell information, där sådan sekretess föreskrivs i nationell lagstiftning eller gemenskapslagstiftning i syfte att skydda legitima ekonomiska intressen, inbegripet det allmänna intresset att behålla sekretess för insynsskydd för statistiska uppgifter och skattesekretess.
...
De skäl till avslag som nämns i [särskilt punkt 2] skall tolkas restriktivt, varvid det i det särskilda fallet skall tas hänsyn till allmänhetens intresse av att informationen lämnas ut. I varje enskilt fall skall allmänhetens intresse av att informationen lämnas ut vägas mot det intresse som betjänas av att begäran avslås. …
...
Miljöinformation som innehas av eller förvaras för offentliga myndigheter och som begärs av en sökande skall tillhandahållas till viss del, där det är möjligt att skilja ut sådana uppgifter som omfattas av punkt 1 d och e eller punkt 2 från den övriga begärda informationen.”
Direktiv 2003/35
I skäl 5 i direktiv 2003/35 anges att unionslagstiftningen bör anpassas till Århuskonventionen med tanke på ratificeringen av konventionen.
Slovakisk rätt
Processrättsliga regler
I artikel 135.1 i civilprocesslagen föreskrivs följande:
… Domstolen är även bunden av avgöranden från Ústavný súd Slovenskej republiky [(den slovakiska författningsdomstolen)] eller från Europeiska domstolen för de mänskliga rättigheterna vilka rör grundläggande rättigheter och friheter.”
I artikel 56.6 i lag nr 38/1993 om inrättande av Ústavný súd Slovenskej republiky samt om dess rättegångsregler och dess domares ställning, i den lydelse som är tillämplig på omständigheterna i det nationella målet, föreskrivs följande:
Om Ústavný súd Slovenskej republiky upphäver ett avgörande eller någon annan giltig åtgärd samt återförvisar målet eller ärendet är den myndighet som har meddelat avgörandet eller vidtagit åtgärden skyldigt att pröva och avgöra målet eller ärendet på nytt. I ett sådant förfarande eller steg är denna myndighet bunden av den právny názor [rättsliga bedömning] som Ústavný súd Slovenskej republiky gjort.”
Bestämmelserna om miljökonsekvensbedömning, stadsplanering och integrerade tillstånd
Lag nr 24/2006
I artikel 1.1 i lag nr 24/2006 om miljökonsekvensbedömning och om ändring av flera lagar, i den lydelse som är tillämplig på omständigheterna i det nationella målet, föreskrivs följande:
Denna lag reglerar
förfarandet för miljökonsekvensbedömning som görs av experter och av allmänheten
...
av planerad verksamhet, innan det beslutas om påbörjande av verksamheten eller innan det beviljas tillstånd för verksamheten i enlighet med särskild lagstiftning.
...”
I artikel 37 i lagen föreskrivs följande:
...
Giltighetstiden för ett slutligt utlåtande avseende en verksamhet är tre år räknat från dess utfärdande. Det slutliga utlåtandet bibehåller sin giltighet om det under denna treårsperiod inleds ett förfarande för påbörjande av eller beviljande av tillstånd för verksamheten i enlighet med särskild lagstiftning.
Giltighetstiden för det slutliga utlåtandet för en verksamhet kan förlängas med en period på två år, vilken kan förnyas på ansökan av sökanden om denne inkommer med skriftlig bevisning för att den planerade verksamheten och de förhållanden som råder på platsen inte har ändrats väsentligt, att det inte har uppkommit några nya fakta som rör det materiella innehållet i miljökonsekvensbeskrivningen av verksamheten och att det inte har utvecklats någon ny teknologi för genomförande av den planerade verksamheten. Beslut om förlängning av giltighetstiden för det slutliga utlåtandet avseende verksamheten ska fattas av det behöriga organet.”
I artikel 65.5 i lagen föreskrivs följande:
Om det slutliga utlåtandet har utfärdats före den 1 februari 2006 och om tillståndsförfarandet för den verksamhet som bedömts inte har inletts i enlighet med den särskilda lagstiftningen härom ska det inges ansökan till ministeriet om förlängning av utlåtandets giltighetstid, i enlighet med vad som anges i artikel 37.7.”
Lag nr 50/1976
I artikel 32 i lag nr 50/1976 om stadsplanering, i den lydelse som är tillämplig på omständigheterna i det nationella målet, föreskrivs följande:
Lokalisering av nybyggnation, ändring av markanvändningen och skyddande av viktiga intressen vad avser markområdet kräver att det har meddelats ett stadsplaneringsbeslut i form av ett
beslut om lokalisering av nybyggnation
...”
Lag nr 245/2003
I artikel 8.3 och 8.4 i lag nr 245/2003 om integrerade åtgärder för förebyggande och bekämpning av miljöföroreningar och om ändring av vissa lagar, i dess lydelse enligt lag nr 532/2005 (nedan kallad lag nr 245/2003), föreskrivs följande:
3)   I de fall då det är fråga om ett integrerat driftstillstånd, vilket förutsätter att det även finns ett tillstånd till uppförande av en nybyggnation eller till ändring av en befintlig byggnation, innefattar förfarandet även ett stadsplaneringsförfarande, ett förfarande för ändringar som företas före byggnationens färdigställande och ett förfarande för tillstånd till inredningsarbeten.
Stadsplaneringsförfarandet, miljökonsekvensbedömningen av anläggningen och fastställandet av villkor till förebyggande av allvarliga industriskador ingår inte i det integrerade tillståndet.”
I artikel 11.2 i lagen föreskrivs följande:
Följande handlingar ska bifogas ansökan [om integrerat tillstånd]:
...
det slutliga utlåtandet i förfarandet för miljökonsekvensbedömning, om driften av den aktuella verksamheten kräver att en sådan bedömning görs,
…
stadsplaneringsbeslutet, om det rör sig om en ny verksamhet eller utbyggnad av en befintlig verksamhet ...”
I artikel 12 i lagen, som har rubriken ”Inledning av förfarandet”, föreskrivs följande:
...
Efter det att det konstaterats att ansökan är fullständig och efter det att parterna i förfarandet och de behöriga organen identifierats ska myndigheten
...
... dels offentliggöra ansökan på dess webbplats, med undantag av de bilagor som inte finns tillgängliga i elektronisk form, dels anslå – under en period om minst 15 dagar – väsentliga uppgifter om ansökan samt om exploatören och verksamheten på myndighetens officiella anslagstavla,
...”
Målet vid den nationella domstolen och tolkningsfrågorna
Det administrativa förfarandet
Mesto Pezinok antog den 26 juni 1997 den allmänna förordningen nr 2/1997 innehållande en detaljplan. I denna detaljplan framgick bland annat lokaliseringen av en avfallsdeponi i en täkt för utvinning av material till tegeltillverkning, vilken kallades Nová jama (den nya täkten).
På grundval av en miljökonsekvensbeskrivning av den planerade lokaliseringen av avfallsdeponin som lades fram av Pezinské tehelne as den 16 december 1998 gjorde miljöministeriet år 1999 en miljökonsekvensbedömning. Miljöministeriet utfärdade ett slutligt utlåtande den 26 juli 1999.
Den 7 augusti 2002 ingav Ekologická skládka en ansökan till den behöriga avdelningen i Mesto Pezinok om ett stadsplaneringsbeslut avseende lokalisering av en avfallsdeponi i Nová jama.
Den 27 mars 2006 förlängde miljöministeriet, på ansökan av Pezinské tehelne as, giltighetstiden för dess slutliga utlåtande från den 26 juli 1999 till den 1 februari 2008.
Genom beslut av den 30 november 2006, i dess lydelse enligt ett beslut från Krajský stavebný úrad v Bratislave (det regionala stadsplaneringskontoret i Bratislava) av den 7 maj 2007, beviljade Mesto Pezinok Ekologická skládkas ansökan om tillstånd för lokalisering av en avfallsdeponi i Nová jama.
Efter det att Ekologická skládka den 25 september 2007 ingett en ansökan om integrerat tillstånd inledde Slovenská inšpekcia životného prostredia, Inšpektorát životného prostredia Bratislava (den slovakiska miljöinspektionen, miljöinspektoratet i Bratislava) (nedan kallat Inšpektorát) ett integrerat förfarande med stöd av lag nr 245/2003, vilken antagits till införlivande av direktiv 96/61. Den 17 oktober 2007 offentliggjorde Inšpektorát, tillsammans med miljöskyddsmyndigheterna, nämnda ansökan, varvid den fastställde en frist på 30 dagar inom vilken allmänheten och de berörda delarna av statsförvaltningen kunde yttra sig över ansökan.
Klagandena i det nationella målet gjorde gällande att Ekologická skládkas ansökan om integrerat tillstånd var ofullständig, eftersom stadsplaneringsbeslutet avseende lokaliseringen av deponin inte hade bifogats, såsom föreskrivs i artikel 11.2 g i lag nr 245/2003, och Inšpektorát vilandeförklarade således det integrerade förfarandet den 26 november 2007 och förelade Ekologická skládka att inkomma med nämnda beslut.
Ekologická skládka gav in beslutet den 27 december 2007, varvid bolaget uppgav att beslutet skulle betraktas som en affärshemlighet. Mot bakgrund härav underlät Inšpektorát att göra beslutet tillgängligt för klagandena i det nationella målet.
Inšpektorát meddelade den 22 januari 2008 Ekologická skládka ett integrerat tillstånd för uppförande av anläggningen ”Pezinok – avfallsdeponi” och för driften av denna anläggning.
Klagandena i det nationella målet överklagade beslutet till Inšpekcia (miljöinspektionen), det vill säga den överordnade miljöskyddsmyndigheten, vilken utgjorde överklagandeinstans i det aktuella ärendet. Inšpekcia beslutade att offentliggöra stadsplaneringsbeslutet om lokaliseringen av deponin på sin officiella anslagstavla under perioden den 14 mars till den 14 april 2008.
I det administrativa förfarandet i andra instans gjorde klagandena i det nationella målet bland annat gällande att Inšpektorát gjort sig skyldigt till felaktig rättstillämpning när det inledde det integrerade förfarandet utan att ha tillgång till stadsplaneringsbeslutet om lokaliseringen av deponin och utan att offentliggöra beslutet när det väl hade getts in av det skälet att det påståtts utgöra en affärshemlighet.
Inšpekcia avslog överklagandet i beslut av den 18 augusti 2008.
Domstolsförfarandet
Klagandena i det nationella målet överklagade beslutet från Inšpekcia av den 18 augusti 2008 till Krajský súd Bratislava, regional förvaltningsdomstol i första instans i Bratislava. Krajský súd Bratislava avslog överklagandet genom dom av den 4 december 2008.
Klagandena i det nationella målet överklagade denna dom till Najvyšší súd Slovenskej republiky (Högsta domstolen i Republiken Slovakien).
Najvyšší súd Slovenskej republiky inhiberade det integrerade tillståndet genom beslut av den 6 april 2009.
Genom dom av den 28 maj 2009 upphävde Najvyšší súd Slovenskej Republiky, med ändring av domen från Krajský súd Bratislava, beslutet från Inšpekcia av den 18 augusti 2008 och beslutet från Inšpektorát av den 22 januari 2008, huvudsakligen med den motiveringen att de behöriga myndigheterna inte hade följt reglerna om den berörda allmänhetens deltagande i det integrerade förfarandet och inte hade gjort en tillräckligt omfattande miljökonsekvensbedömning av anläggandet av deponin.
Ekologická skládka väckte talan mot beslutet av den 6 april 2009 och mot domen av den 28 maj 2009 vid Ústavný súd Slovenskej republiky (Republiken Slovakiens författningsdomstol) den 25 juni 2009 respektive den 3 september 2009.
Ústavný súd Slovenskej republiky fann, i dom av den 27 maj 2010, att Najvyšší súd Slovenskej republiky hade åsidosatt Ekologická skládkas grundläggande rätt till domstolsskydd enligt artikel 46.1 i Republiken Slovakiens konstitution, dess grundläggande äganderätt enligt artikel 20.1 i konstitutionen och dess rätt att ostört få nyttja sin egendom enligt artikel 1 i tilläggsprotokollet till Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna, som undertecknades i Rom den 4 november 1950.
Ústavný súd Slovenskej republiky ansåg särskilt att Najvyšší súd Slovenskej republiky inte hade beaktat alla principer som gäller för det administrativa förfarandet och att den hade överskridit sina befogenheter när den prövade lagenligheten av förfarandet och av beslutet om miljökonsekvensbedömning trots att klagandena inte hade bestritt denna och att den inte hade någon behörighet att uttala sig i denna fråga.
I sin dom upphävde Ústavný súd Slovenskej republiky således det angripna beslutet och den angripna domen samt återförvisade målet till Najvyšší súd Slovenskej republiky för ny prövning.
Enligt Najvyšší súd Slovenskej republiky anser flera deltagare i rättegången i det nationella målet att den är bunden av domen från Ústavný súd Slovenskej republiky av den 27 maj 2010. Najvyšší súd Slovenskej republiky har emellertid angett att den fortfarande hyser tvivel om huruvida de angripna avgörandena är förenliga med unionsrätten.
Mot denna bakgrund beslutade Najvyšší súd Slovenskej republiky att vilandeförklara målet och att ställa följande frågor till domstolen:
1)
Innebär [unions]rätten (närmare bestämt artikel 267 FEUF) en skyldighet eller en rättighet för högsta domstolen i en medlemsstat att ’på eget initiativ’ begära förhandsavgörande från [EU-domstolen] även i ett skede i domstolsförfarandet då författningsdomstolen har upphävt en dom av högsta domstolen, som huvudsakligen grundas på tillämpningen av [unionsrätten] på miljöskyddsområdet, och ålagt högsta domstolen att följa författningsdomstolens bedömning att de rättigheter, såväl processuella som materiella, som enligt författningen tillkommer en deltagare i rättegången har åsidosatts, utan att författningsdomstolen tagit hänsyn till de [unionsrättsliga] aspekterna i målet, det vill säga då författningsdomstolen som högsta rättsinstans inte har funnit det nödvändigt att begära förhandsavgörande från [EU-domstolen] och på förhand har uteslutit att rätten till en god miljö och skyddet härför gör sig gällande i målet?
Är det möjligt att uppnå det grundläggande syftet med de samordnade åtgärderna för förebyggande som särskilt föreskrivs i skälen 8, 9 och 23 i ingressen till … direktiv [96/61] och i artiklarna 1 och 15 i direktivet samt generellt i [unionsrätten] på miljöområdet – det vill säga förebyggande och bekämpning av föroreningar även med hjälp av allmänhetens deltagande i förverkligandet av en hög skyddsnivå för miljön som helhet – när den berörda allmänheten inte vid tiden för inledandet av förfarandet för samordnat förebyggande har tillgång till alla relevanta handlingar (artikel 6 jämförd med artikel 15 i direktiv [96/61]), däribland särskilt beslutet om lokaliseringen av en anläggning (avfallsdeponi), men när sökanden senare under förfarandet i första instans bifogar den handling som saknas på villkoret att den inte lämnas ut till övriga parter i förfarandet, eftersom det är fråga om en affärshemlighet, trots att det rimligen kan antas att beslutet om lokalisering av anläggningen (och särskilt skälen för beslutet) skulle ha en väsentlig inverkan på de förslag, synpunkter och andra kommentarer som kan komma att lämnas?
Uppfylls målen med … direktiv [85/337] – särskilt med beaktande av [unionsrätten] på miljöområdet, närmare bestämt kravet i artikel 2 i direktivet att projekt ska bli föremål för en bedömning av deras miljöpåverkan innan tillstånd meddelas – i en situation där ett ursprungligt utlåtande från miljöministeriet, vilket utfärdades år 1999 och avslutade förfarandet för miljökonsekvensbedömning, förlängs flera år senare genom ett beslut utan att en ny miljökonsekvensbedömning görs? Uttryckt på ett annat sätt, kan det antas att ett beslut som har fattats i enlighet med direktiv [85/337] har obegränsad giltighet?
Är det generella kravet, som föreskrivs i direktiv [96/61] (särskilt i ingressen och i artiklarna 1 och 15a) – enligt vilket varje medlemsstat ska säkerställa förebyggande och bekämpning av föroreningar även genom att ge den berörda allmänheten möjlighet att i rimlig tid använda sig av ett rättvist och opartiskt administrativt rättsmedel samt att få till stånd en rättvis och opartisk domstolsprövning – i förening med artikel 10a i direktiv [85/337] och artiklarna 6 samt 9.2 och 9.4 i Århuskonventionen, tillämpligt på allmänhetens möjlighet att hos förvaltningsmyndighet eller domstol begära interimistiska åtgärder i enlighet med nationell rätt (exempelvis ett beslut om inhibition av ett samordnat tillstånd) som gör det möjligt att interimistiskt, det vill säga fram till dess att saken slutligt avgörs, ställa in genomförandet av den verksamhet som tillståndsansökan avser?
Är det möjligt att ett domstolsavgörande, som uppfyller kraven i direktiv [96/61], direktiv [85/337] eller artikel 9.2–9.4 i Århuskonventionen när det gäller allmänhetens rätt enligt dessa bestämmelser till ett rättvist domstolsskydd i den mening som avses i artikel 191.1 och 191.2 [FEUF] avseende Europeiska unionens miljöpolitik, samtidigt kan innebära en otillåten kränkning av exploatörens äganderätt till en anläggning, såsom den bland annat säkerställs i artikel 1 i tilläggsprotokollet till Europeiska konventionen om mänskliga rättigheter och grundläggande friheter, till exempel genom att ett giltigt integrerat tillstånd till driften av en ny anläggning som en sökande beviljats upphävs i domstolsförfarandet?”
Prövning av tolkningsfrågorna
Upptagande till sakprövning
Inšpekcia, Ekologická skládka och den slovakiska regeringen har, på olika grunder, hävdat att begäran om förhandsavgörande eller vissa av de frågor som ställts inte kan prövas i sak.
Enligt Inšpekcia och Ekologická skládka ska begäran om förhandsavgörande avvisas i sin helhet, eftersom alla tolkningsfrågorna avser situationer som i samtliga delar regleras av nationell rätt, särskilt av de rättsakter som antagits till införlivande av direktiven 85/337 och 96/61. Enligt Ekologická skládka följer det härav att dessa direktiv saknar direkt effekt, medan Inšpekcia anser att direktiven är tillräckligt klara för att begäran om förhandsavgörande ska anses obehövlig. Inšpekcia har även hävdat att tolkningsfrågorna skulle ha ställts i det inledande skedet i förfarandet vid Najvyšší súd Slovenskej republiky. Ekologická skládka anser likaledes att frågorna är överflödiga, eftersom Najvyšší súd Slovenskej republiky ändå är bunden av den ståndpunkt som Ústavný súd Slovenskej republiky intagit och eftersom ingen av parterna i det nationella målet har anmodat om att frågorna ska hänskjutas till EU-domstolen för förhandsavgörande.
Ekologická skládka har vidare gjort gällande att den åtskillnad som görs i nationell rätt mellan det integrerade förfarandet, stadsplaneringsförfarandet och miljökonsekvensbedömningen innebär att den andra och den tredje frågan saknar relevans för avgörandet av det nationella målet. Enligt Inšpekcia utgör denna åtskillnad grund för att avvisa den tredje, den fjärde och den femte frågan. Den innebär nämligen att ett fel eller en brist i stadsplaneringsbeslutet eller i miljökonsekvensbedömningen inte påverkar lagenligheten av det integrerade tillståndet.
Härutöver anser Ekologická skládka och den slovakiska regeringen att den fjärde frågan är hypotetisk. De interimistiska åtgärder som Najvyšší súd Slovenskej republiky har förordnat om i sitt beslut av den 6 april 2009 har helt förlorat sin verkan. Dessutom saknar frågan relevans i det mål som den hänskjutande domstolen har att avgöra, eftersom det nationella målet inte avser förordnande om nya interimistiska åtgärder, utan snarare giltigheten av de angripna förvaltningsbesluten.
Ekologická skládka har slutligen hävdat att även den femte frågan är hypotetisk, eftersom den avser det avgörande som Najvyšší súd Slovenskej republiky har att fatta då det nationella målet ska avgöras i sak. Dessutom ska denna fråga även avvisas av det skälet att den avser tolkningen av nationell konstitutionell rätt.
I detta hänseende ska det erinras om att det enligt fast rättspraxis uteslutande ankommer på den nationella domstolen, vid vilken tvisten anhängiggjorts och vilken har ansvaret för det rättsliga avgörandet, att mot bakgrund av de särskilda omständigheterna i målet bedöma såväl om ett förhandsavgörande är nödvändigt för att döma i saken som relevansen av de frågor som ställs till domstolen. Domstolen är följaktligen i princip skyldig att meddela ett förhandsavgörande när de frågor som ställts av den nationella domstolen avser tolkningen av unionsrätten (dom av den 10 mars 2009 i mål C-169/07, Hartlauer, REG 2009, s. I-1721, punkt 24, och av den 19 juli 2012 i mål C-470/11, Garkalns, punkt 17).
Frågor om tolkningen av unionsrätten presumeras således vara relevanta. En tolkningsfråga från en nationell domstol kan enbart avvisas då det är uppenbart att den begärda tolkningen av unionsrätten inte har något samband med de verkliga omständigheterna eller föremålet för tvisten vid den nationella domstolen eller då frågorna är hypotetiska eller EU-domstolen inte har tillgång till sådana uppgifter om de faktiska eller rättsliga omständigheterna som är nödvändiga för att kunna ge ett användbart svar på de frågor som ställts till den (dom av den 1 juni 2010 i de förenade målen C-570/07 och C-571/07, Blanco Pérez och Chao Gómez, REU 2010, s. I-4629, punkt 36, och av den 5 juli 2012 i mål C-509/10, Geistbeck, punkt 48).
Argumentet att den aktuella frågan regleras fullt ut i nationell rätt kan emellertid inte läggas till grund för slutsatsen att det är uppenbart att tolkningen av de unionsrättsliga regler som nämnts av den nationella domstolen inte har något samband med tvisten vid den nationella domstolen. Detta gör sig än mer gällande eftersom det är utrett att de tillämpliga nationella bestämmelserna till viss del har antagits till införlivande av unionsrättsakter. Detta argument kan således inte motbevisa den presumtion avseende relevans som har nämnts i föregående punkt.
Det kan vidare konstateras att det faktum att de aktuella direktiven, enligt vad som påståtts, saknar direkt effekt inte påverkar denna analys, eftersom domstolen enligt artikel 267 FEUF är behörig att döma i frågor om förhandsavgörande avseende tolkningen av rättsakter som antagits av unionens institutioner, oavsett om de är direkt tillämpliga eller inte (dom av den 10 juli 1997 i mål C-373/95, Maso m.fl., REG 1997, s. I-4051, punkt 28, av den 16 juli 2009 i mål C-254/08, Futura Immobiliare m.fl., REG 2009, s. I-6995, punkt 34, och av den 27 november 2012 i mål C-370/12, Pringle, punkt 89). När det vidare gäller påståendet att de tillämpliga reglerna är klara och att det därför inte är ändamålsenligt att begära förhandsavgörande, ska det erinras om att artikel 267 FEUF alltid tillåter en nationell domstol – om denna anser det lämpligt – att hänskjuta tolkningsfrågor till EU-domstolen (se, för ett liknande resonemang, dom av den 26 maj 2011 i de förenade målen C-165/09–C-167/09, Stichting Natuur en Milieu m.fl., REU 2011, s. I-4599, punkt 52 och där angiven rättspraxis).
Övriga argument som Inšpekcia och Ekologická skládka anfört till stöd för att begäran om förhandsavgörande ska avvisas i sin helhet avser föremålet för den första frågan och kommer att behandlas i samband med att domstolen prövar denna fråga.
När det gäller det faktum att det görs åtskillnad mellan olika förfaranden i nationell rätt ska det noteras att den nationella domstolen har en helt annan uppfattning om konsekvenserna härav än Inšpekcia och Ekologická skládka. I förfaranden enligt artikel 267 FEUF råder emellertid tydlig åtskillnad mellan EU-domstolens och den nationella domstolens funktioner och den sistnämnda är ensam behörig att tolka den nationella lagstiftningen (dom av den 17 juni 1999 i mål C-295/97, Piaggio, REG 1999, s. I-3735, punkt 29, och av den 17 juli 2008 i mål C-500/06, Corporación Dermoestética, REG 2008, s. I-5785, punkt 21). Nämnda faktum innebär således inte i sig att det måste anses uppenbart att de ställda frågorna saknar samband med de verkliga omständigheterna eller föremålet för den aktuella tvisten.
Vad gäller huruvida den fjärde frågan kan prövas framgår det av beslutet om hänskjutande att Najvyšší súd Slovenskej republiky har förordnat om nya interimistiska åtgärder innebärande inhibition av de beslut som det nationella målet rör. Ekologická skládka har dessutom angett i sitt skriftliga yttrande att den fann det nödvändigt att väcka talan mot nämna åtgärder. Mot bakgrund härav kan den fjärde frågan inte anses vara hypotetisk.
När det slutligen gäller frågan huruvida den femte frågan kan prövas är det utrett att Ústavný súd Slovenskej republiky fann att Najvyšší súd Slovenskej republiky hade åsidosatt Ekologická skládkas äganderätt genom sin dom av den 28 maj 2009, varigenom det konstaterades att det integrerade tillståndet hade beviljats på ett sätt som inte var förenligt med unionsrätten. Eftersom den nationella domstolen fortfarande hyser tvivel om huruvida de i det nationella målet angripna besluten är förenliga med unionsrätten kan den femte frågan inte anses vara rent hypotetisk. Dessutom framgår det av lydelsen av denna fråga att den inte avser tolkning av nationell konstitutionell rätt.
De frågor som den nationella domstolen har ställt kan således prövas i sak.
Den första frågan
Najvyšší súd Slovenskej republiky har ställt den första frågan för att få klarhet i huruvida artikel 267 FEUF ska tolkas så, att en nationell domstol på eget initiativ kan begära förhandsavgörande från EU-domstolen även om det mål den har att avgöra har återförvisats till den efter det att dess första avgörande i saken upphävts av författningsdomstolen i den aktuella medlemsstaten och den, enligt en nationell bestämmelse, är skyldig att lägga författningsdomstolens rättsliga bedömning till grund för sitt avgörande av tvisten. Najvyšší súd Slovenskej republiky önskar även få klarhet i huruvida artikel 267 FEUF ska tolkas så, att en sådan nationell domstol är skyldig att begära förhandsavgörande från EU-domstolen fastän dess avgöranden kan bli föremål för en talan vid en författningsdomstol, vilken är begränsad till prövningen av om de rättigheter och friheter som följer av den nationella konstitutionen eller av en internationell konvention har åsidosatts.
Inledningsvis finner domstolen att Najvyšší súd Slovenskej republiky, genom sin första fråga, även önskar få klarhet i huruvida den enligt unionsrätten kan underlåta att tillämpa en nationell bestämmelse enligt vilken den inte får beakta en grund avseende åsidosättande av unionsrätten som inte har åberopats av parterna i det nationella målet. Det framgår emellertid av beslutet om hänskjutande att denna frågeställning endast avser direktiv 85/337 och således endast ska besvaras om det, med hänsyn till svaret på den tredje frågan, visar sig att detta direktiv är tillämpligt i det nationella målet.
När det gäller övriga aspekter av den första tolkningsfrågan framgår det av rättspraxis att en nationell domstol enligt artikel 267 FEUF har en mycket vittgående möjlighet att hänskjuta en fråga till EU-domstolen, om den bedömer att det i ett mål som pågår inför den har uppkommit frågor som kräver ett avgörande avseende tolkningen eller giltigheten av bestämmelser i unionsrätten för att den ska kunna döma i målet (dom av den 27 juni 1991 i mål C-348/89, Mecanarte, REG 1991, s. I-3277, punkt 44, och av den 5 oktober 2010 i mål C-173/09, Elchinov, REU 2010, s. I-8889, punkt 26).
Artikel 267 FEUF ger således en nationell domstol en möjlighet, och i förekommande fall en skyldighet, att begära förhandsavgörande så snart den, antingen på eget initiativ eller på begäran av parterna i målet, finner att saken i målet rör en fråga som avses i första stycket i denna artikel (dom av den 10 juli 1997 i mål C-261/95, Palmisani, REG 1995, s. I-4025, punkt 20, och av den 21 juli 2011 i mål C-104/10, Kelly, REU 2011, s. I-6813, punkt 61). Därmed hindrar den omständigheten att parterna i det nationella målet inte har väckt någon unionsrättslig fråga inför den nationella domstolen inte att det begärs förhandsavgörande från EU-domstolen (dom av den 16 juni 1981 i mål 126/80, Salonia, REG 1981, s. 1563, punkt 7, svensk specialutgåva, volym 6, s. 129, och av den 8 mars 2012 i mål C-251/11, Huet, punkt 23).
Begäran om förhandsavgörande vilar nämligen på en dialog mellan domstolar. Denna dialog kommer endast till stånd om den nationella domstolen finner att det är relevant och nödvändigt att framställa en sådan begäran (dom av den 16 december 2008 i mål C-210/06, Cartesio, REG 2008, s. I-9641, punkt 91, och av den 9 november 2010 i mål C-137/08, VB Pénzügyi Lízing, REU 2010, s. I-10847, punkt 29).
Dessutom kan förekomsten av en nationell processrättslig regel inte påverka möjligheten för en nationell domstol att begära förhandsavgörande från EU-domstolen när den, såsom i det nationella målet, är osäker på hur unionsrätten ska tolkas (domen i det ovannämnda målet Elchinov, punkt 25, och av den 20 oktober 2011 i mål C-396/09, Interedil, REU 2011, s. I-9915, punkt 35).
En nationell bestämmelse, enligt vilken en domstol är bunden av en högre instans rättsliga bedömning, hindrar således inte den förstnämnda domstolen från att till EU-domstolen ställa frågor om tolkningen av de delar av unionsrätten som den rättsliga bedömningen avser. Det måste nämligen stå en sådan domstol fritt att ställa frågor till EU-domstolen, om den anser att ett avgörande i enlighet med den högre instansen rättsliga bedömning skulle strida mot unionsrätten (dom av den 9 mars 2010 i mål C-378/08, ERG m.fl., REU 2010, s. I-1919, punkt 32, samt domen i det ovannämnda målet Elchinov, punkt 27).
En nationell domstol som har utnyttjat sin möjlighet enligt artikel 267 FEUF är bunden av EU-domstolens tolkning av de aktuella bestämmelserna när den avgör tvisten i det mål som är anhängigt vid den och är, i förekommande fall, skyldig att avvika från den högre instansens bedömning om den mot bakgrund av EU-domstolens tolkning finner att denna bedömning är oförenlig med unionsrätten (domen i det ovannämnda målet Elchinov, punkt 30).
De principer som nämnts i de föregående punkterna gör sig även gällande för Najvyšší súd Slovenskej republiky vad gäller den rättsliga bedömning som författningsdomstolen i den aktuella medlemsstaten gjort i det nationella målet. Enligt fast rättspraxis får nämligen bestämmelser i nationell rätt inte, ens om de har rang av grundlag, undergräva unionsrättens enhetlighet och effektivitet (dom av den 17 december 1970 i mål 11/70, Internationale Handelsgesellschaft, REG 1970, s. 1125, punkt 3, svensk specialutgåva, volym 1, s. 503, och av den 8 september 2010 i mål C-409/06, Winner Wetten, REU 2010, s. I-8015, punkt 61). Domstolen har dessutom redan slagit fast att nämnda principer är tillämpliga i förhållandet mellan en författningsdomstol och övriga nationella domstolar (dom av den 22 juni 2010 i de förenade målen C-188/10 och C-189/10, Melki och Abdeli, REU 2010, s. I-5667, punkterna 41–45).
Den nationella bestämmelse enligt vilken Najvyšší súd Slovenskej republiky är skyldig att rätta sig efter Ústavný súd Slovenskej republikys rättsliga bedömning kan således inte hindra förstnämnda domstol från att, närhelst under förfarandet den finner det lämpligt, begära förhandsavgörande från EU-domstolen och att, i förekommande fall, avvika från Ústavný súd Slovenskej republikys bedömning i den mån som den anser den strida mot unionsrätten.
Najvyšší súd Slovenskej republiky är, i egenskap av högsta domstolsinstans, till och med skyldig att begära förhandsavgörande från EU-domstolen så snart den finner att saken i målet rör en fråga som avses i första stycket i artikel 267 FEUF. Möjligheten att väcka talan vid författningsdomstolen i den aktuella medlemsstaten mot ett avgörande från en nationell domstol, varvid författningsdomstolen endast kan pröva om de rättigheter och friheter som följer av den nationella konstitutionen eller av en internationell konvention har åsidosatts, innebär nämligen inte att den nationella domstolen inte kan kvalificeras som en domstol mot vars avgöranden det inte finns något rättsmedel enligt nationell lagstiftning i den mening som avses i artikel 267 tredje stycket FEUF.
Mot denna bakgrund ska den första frågan besvaras enligt följande: Artikel 267 FEUF ska tolkas så, att en nationell domstol, såsom den hänskjutande domstolen, är skyldig att på eget initiativ begära förhandsavgörande från EU-domstolen trots att det mål den har att avgöra har återförvisats till den efter det att dess första avgörande i saken upphävts av författningsdomstolen i den aktuella medlemsstaten och trots att den, enligt en nationell bestämmelse, är skyldig att lägga författningsdomstolens rättsliga bedömning till grund för sitt avgörande av tvisten.
Den andra frågan
Den nationella domstolen har ställt den andra frågan för att få klarhet i huruvida direktiv 96/91 ska tolkas så, att det kräver att den berörda allmänheten, redan från det att tillståndsförfarandet avseende en deponi inleds, ges tillgång till ett stadsplaneringsbeslut om lokalisering av anläggningen. Den vill även få klarhet i huruvida en vägran att tillhandahålla detta beslut kan vara motiverad av det skälet att informationen i beslutet påstås omfattas av skyddet för affärshemligheter eller, om så inte är fallet, huruvida den felaktighet som begåtts kan rättas till genom att den berörda allmänheten ges möjlighet att ta del av beslutet under det administrativa förfarandet i andra instans.
Inledningsvis kan det konstateras att det framgår av beslutet om hänskjutande att den anläggning som det nationella målet avser är en deponi som dagligen mottar mer än 10 ton avfall och som har en samlad kapacitet på över 25000 ton avfall. Den omfattas således av tillämpningsområdet för direktiv 96/61, såsom detta framgår av artikel 1 i direktivet i förening med punkt 5.4 i bilaga 1 till direktivet.
I artikel 15 i direktiv 96/61 föreskrivs att den berörda allmänheten ska ges tillfälle att delta i förfaranden för meddelande av tillstånd för nya anläggningar och att villkoren för deltagandet framgår av bilaga V till direktivet. Enligt denna bilaga ska allmänheten upplysas om från vilka myndigheter de kan erhålla relevant information och om när och var denna information kommer att göras tillgänglig.
Dessa bestämmelser om allmänhetens deltagande ska tolkas mot bakgrund av – och med beaktande av – bestämmelserna i Århuskonventionen, till vilken unionslagstiftningen bör ”anpassas” enligt skäl 5 i direktiv 2003/35, vilket direktiv delvis ändrade direktiv 96/61 (dom av den 12 maj 2011 i mål C-115/09, Bund für Umwelt und Naturschutz Deutschland, Landesverband Nordrhein-Westfalen, REU 2011, s. I-3673, punkt 41). I artikel 6.6 i Århuskonventionen föreskrivs emellertid att allmänheten måste kunna ta del av all information som är av betydelse för beslutsprocessen för tillstånd till sådan verksamhet som avses i bilaga I till konventionen, såsom exempelvis deponier som tar emot mer än 10 ton avfall per dygn eller med en total kapacitet som överstiger 25000 ton avfall.
Den allmänhet som berörs av det tillståndsförfarande som avses i direktiv 96/91 måste, i princip, kunna få tillgång till alla uppgifter som är relevanta för förfarandet.
Det framgår av beslutet om hänskjutande och av de handlingar som getts in till domstolen att stadsplaneringsbeslutet om lokalisering av den anläggning som det nationella målet avser ingår i underlaget för det slutliga beslutet att tillåta eller inte tillåta att anläggningen uppförs och att detta beslut innehåller uppgifter om den planerade anläggningens inverkan på miljön, om de villkor som exploatören ålagts att följa för att begränsa denna inverkan, om de invändningar som parterna i stadsplaneringsförfarandet framfört och om skälen till de val den behöriga myndigheten träffat vid antagandet av beslutet. Dessutom krävs det enligt de tillämpliga nationella bestämmelserna att stadsplaneringsbeslutet bifogas den tillståndsansökan som skickas till den behöriga myndigheten. Härav följer att beslutet måste anses innehålla relevant information i den mening som avses i bilaga V till direktiv 96/61 och att den berörda allmänheten således i princip måste kunna få tillgång till det under tillståndsförfarandet för nämnda anläggning.
Det framgår av artikel 15.4 i direktiv 96/61 att den berörda allmänhetens deltagande kan inskränkas genom de begränsningar som föreskrivs i artikel 3.2 och 3.3 i direktiv 90/313. Vid tidpunkten för omständigheterna i det nationella målet hade direktiv 90/313 emellertid upphävts och ersatts av direktiv 2003/4. Med beaktande av den jämförelsetabell som bifogats direktiv 2003/4, skyldigheten att anpassa unionslagstiftningen till Århuskonventionen och den utformning artikel 15 i direktiv 96/61 fick vid den senaste kodifieringen genom Europaparlamentets och rådets direktiv 2008/1/EG av den 15 januari 2008 om samordnade åtgärder för att förebygga och begränsa föroreningar (EUT L 24, s. 8) måste artikel 15.4 i direktiv 96/61 tolkas så, att den hänvisar till de begränsningar som föreskrivs i artikel 4.1, 4.2 och 4.4 i direktiv 2003/4.
Enligt artikel 4.2 första stycket d i direktiv 2003/4 får medlemsstaterna föreskriva att begäran om miljöinformation ska avslås, om utlämnande av informationen skulle ha negativa följder för sekretess som omfattar kommersiell eller industriell information, där sådan sekretess föreskrivs i nationell lagstiftning eller unionslagstiftning i syfte att skydda legitima ekonomiska intressen.
Med hänsyn bland annat till att lokalisering av de verksamheter som avses i direktiv 96/91 är av stor vikt, och såsom framgår av punkt 79 i denna dom, är så emellertid inte fallet när det gäller ett beslut genom vilket en myndighet beviljar tillstånd, utifrån tillämpliga bestämmelser om stadsplanering, till lokalisering av en anläggning som omfattas av tillämpningsområdet för detta direktiv.
Även om det skulle antas att vissa delar av skälen till ett stadsplaneringsbeslut i undantagsfall skulle kunna innehålla kommersiell eller industriell information som omfattas av sekretess är det i förevarande fall utrett att sekretesskyddet för sådana uppgifter har åberopats som grund för att inte ge den berörda allmänheten tillgång till någon del över huvud taget av stadsplaneringsbeslutet om lokalisering av den anläggning som det nationella målet avser, vilket strider mot artikel 4.4 i direktiv 2003/4.
Härav följer att det faktum att stadsplaneringsbeslutet om lokalisering av den anläggning som det nationella målet avser inte gjordes tillgängligt för den berörda allmänheten under det administrativa förfarandet i första instans inte kunde motiveras med hänvisning till undantaget i artikel 15.4 i direktiv 96/61. Det är således nödvändigt för Najvyšší súd Slovenskej republiky att få klarhet i huruvida detta fel i det administrativa förfarandet i första instans kunde rättas till genom att den berörda allmänheten fick möjlighet att ta del av beslutet under det administrativa förfarandet i andra instans och huruvida ett åsidosättande av artikel 15 i direktiv 96/94 därmed kunde undvikas.
I avsaknad av gemenskapsbestämmelser/unionsbestämmelser på området ankommer det på varje medlemsstat att i sin rättsordning fastställa de processuella regler som gäller för talan i domstol och andra förfaranden som syftar till att säkerställa skyddet av de rättigheter för enskilda som följer av unionsrätten. Dessa regler får emellertid varken vara mindre förmånliga än de som avser liknande talan som grundas på nationell rätt (likvärdighetsprincipen) eller medföra att det i praktiken blir omöjligt eller orimligt svårt att utöva rättigheter som följer av unionsrätten (effektivitetsprincipen) (dom av den 14 december 1995 i mål C-312/93, Peterbroeck, REG 1995, s. I-4599, punkt 12, och av den 12 juli 2012 i mål C-378/10, VALE Építési, punkt 48 och där angiven rättspraxis).
Enligt likvärdighetsprincipen krävs att alla regler avseende talan i domstol eller andra förfaranden ska tillämpas på samma sätt oavsett om talan respektive ansökan grundar sig på åsidosättande av unionsrätten eller på åsidosättande av nationell rätt (se, bland annat, dom av 19 juli 2012 i mål C-591/10, Littlewoods Retail m.fl., punkt 31, och av den 4 oktober 2012 i mål C-249/11, Byankov, punkt 70). Det ankommer således på den nationella domstolen att pröva huruvida det enligt nationell rätt är möjligt att rätta till jämförbara förfarandefel, som innebär avvikelse från nationell rätt, under det administrativa förfarandet i andra instans.
Även om unionsrätten inte utgör hinder för att det enligt nationella bestämmelser i vissa fall kan vara tillåtet att i efterhand rätta till åtgärder eller handlingar som strider mot unionsrätten är en sådan möjlighet villkorad av att den inte möjliggör för de berörda att kringgå de unionsrättsliga bestämmelserna eller att undgå deras tillämpning och att denna möjlighet förblir ett undantag (dom av den 3 juli 2008 i mål C-215/06, kommissionen mot Irland, REG 2008, s. I-4911, punkt 57).
Enligt artikel 15 i direktiv 96/61 ska medlemsstaterna se till att den berörda allmänheten på ett tidigt stadium ges tillfälle att på ett effektivt sätt delta i tillståndsförfarandet. Denna bestämmelse ska tolkas mot bakgrund av skäl 23 i direktivet, enligt vilken allmänheten bör ges tillgång till information som rör tillståndsansökningar rörande nya anläggningar innan det fattas beslut härom och artikel 6 i Århuskonventionen. Enligt sistnämnda artikel ska deltagandet ske på ett tidigt stadium, det vill säga när alla alternativ är möjliga och allmänheten kan delta på ett meningsfullt sätt, och allmänheten ska ges tillgång till all information som är av betydelse så snart den blir tillgänglig. Härav följer att den berörda allmänheten ska kunna ta del av alla relevanta uppgifter redan i det administrativa förfarandet i första instans och innan det första beslutet antas, såvitt dessa uppgifter är tillgängliga i detta skede i förfarandet.
När det gäller frågan huruvida effektivitetsprincipen utgör hinder för att ett fel rättas till under förfarandet i andra instans genom att allmänheten ges möjlighet att ta del av relevanta handlingar som inte var tillgängliga under det administrativa förfarandet i första instans, framgår det av de uppgifter som lämnats av Najvyšší súd Slovenskej republiky att förvaltningsmyndigheten i andra instans, enligt den tillämpliga nationella lagstiftningen, har behörighet att ändra det förvaltningsbeslut som meddelats i första instans. Det ankommer emellertid på Najvyšší súd Slovenskej republiky att pröva huruvida alla alternativ fortfarande är möjliga, i den mening som avses i artikel 15.1 i direktiv 96/91 tolkad mot bakgrund av artikel 6.4 i Århuskonventionen, under det administrativa förfarandet i andra instans. Najvyšší súd Slovenskej republiky har även att pröva huruvida en rättelse i detta skede av förfarandet, genom att den berörda allmänheten ges möjlighet att ta del av relevanta handlingar, innebär att allmänheten fortfarande kan delta på ett meningsfullt sätt i beslutsförfarandet.
Effektivitetsprincipen utgör följaktligen inte hinder för att en oberättigad vägran att ge den berörda allmänheten tillgång till det stadsplaneringsbeslut som det nationella målet avser under det administrativa förfarandet i första instans kan rättas till under det administrativa förfarandet i andra instans, under förutsättning att alla alternativ fortfarande är möjliga och att en rättelse i detta skede i förfarandet innebär att allmänheten fortfarande kan delta på ett meningsfullt sätt i beslutsförfarandet. Det ankommer på den nationella domstolen att pröva huruvida så är fallet.
Mot denna bakgrund ska den andra frågan besvaras enligt följande: Direktiv 96/61 ska tolkas så, att det
kräver att den berörda allmänheten ges tillgång till ett stadsplaneringsbeslut, såsom det som är i fråga i det nationella målet, redan från det att tillståndsförfarandet avseende den aktuella anläggningen inleds,
inte tillåter att de behöriga nationella myndigheterna nekar den berörda allmänheten tillgång till ett sådant beslut med hänvisning till skyddet för sekretess som omfattar kommersiell eller industriell information, där sådan sekretess föreskrivs i nationell lagstiftning eller unionslagstiftning i syfte att skydda legitima ekonomiska intressen, och
inte utgör hinder för att en oberättigad vägran att ge den berörda allmänheten tillgång till ett sådant stadsplaneringsbeslut som det nationella målet avser under det administrativa förfarandet i första instans, kan rättas till under det administrativa förfarandet i andra instans, under förutsättning att alla alternativ fortfarande är möjliga och att en rättelse i detta skede i förfarandet innebär att allmänheten fortfarande kan delta på ett meningsfullt sätt i beslutsförfarandet. Det ankommer på den nationella domstolen att pröva huruvida så är fallet.
Den tredje frågan
Den nationella domstolen har ställt den tredje frågan för att få klarhet i huruvida direktiv 85/337 ska tolkas så, att det utgör hinder för att giltighetstiden för ett utlåtande inom ramen för en miljökonsekvensbedömning av ett projekt på ett giltigt sätt kan förlängas flera år efter det att det utfärdades och huruvida det enligt direktivet krävs att det i så fall görs en ny miljökonsekvensbedömning av projektet.
Inšpekcia, liksom den slovakiska och den tjeckiska regeringen, har hävdat att direktiv 85/337 inte är tillämpligt i tidsmässigt hänseende på den situation som avses i det nationella målet.
Enligt fast rättspraxis är principen att projekt som kan antas medföra en betydande miljöpåverkan ska bli föremål för en miljökonsekvensbedömning inte tillämplig när en formell ansökan om tillstånd för ett projekt har getts in innan det att fristen för införlivande av direktiv 85/337 löpt ut (dom av den 11 augusti 1995 i mål C-431/92, kommissionen mot Tyskland, REG 1995, s. I-2189, punkterna 29 och 32, och dom av den 18 juni 1998 i mål C-81/96, Gedeputeerde Staten van Noord-Holland, REG 1998, s. I-3923, punkt 23).
Detta direktiv avser nämligen i stor utsträckning projekt av viss omfattning som ofta tar lång tid att genomföra. Det vore således inte lämpligt att redan komplicerade nationella förfaranden skulle belastas och försenas av särskilda krav i direktivet och att situationer som redan föreligger skulle beröras av detta (se domen i det ovannämnda målet Gedeputeerde Staten van Noord Holland, punkt 24).
I förevarande fall framgår det av de handlingar som getts in till domstolen att exploatörens första åtgärd för att utverka tillstånd till genomförande av projektet avseende den deponi som det nationella målet avser vidtogs den 16 december 1998 och bestod i ingivandet av en ansökan om en miljökonsekvensbedömning av projektet. Det framgår emellertid av artikel 2 i akten om villkoren för Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens anslutning till de fördrag som ligger till grund för Europeiska unionen och om anpassning av fördragen (EUT L 236, 2003, s. 33) att direktiv 85/337 skulle införlivas av Republiken Slovakien från och med dagen för denna medlemsstats anslutning till unionen, det vill säga den 1 maj 2004.
Det ska emellertid noteras att den slovakiska administrationens beviljande av tillstånd för anläggandet av den deponi som det nationella målet avser har erfordrat tre successiva förfaranden, vilka vart och ett avslutades med att ett beslut antogs.
När det gäller de två första förfarandena inkom exploatörens ansökningar den 16 december 1998 respektive den 7 augusti 2002, det vill säga innan det att fristen för införlivande av direktiv 85/337 hade löpt ut. Ansökan om integrerat tillstånd ingavs däremot inte förrän den 25 september 2007, det vill säga efter utgången av denna frist. Det ska således bedömas huruvida ingivandet av de två första ansökningarna kan anses innebära att tillståndsförfarandet formellt sett inleddes i den mening som avses i den rättspraxis som nämnts i punkt 94 i denna dom.
De ansökningar som getts in under de två första etapperna i förfarandet ska inte förväxlas med informella kontakter, vilka inte innebär att tillståndsförfarandet formellt sett har inletts (se, för ett liknande resonemang, domen i det ovannämnda målet kommissionen mot Tyskland, punkt 32).
Den miljökonsekvensbedömning som avslutades år 1999 gjordes dessutom för att möjliggöra genomförandet av deponiprojektet, vilket var föremål för det integrerade tillståndet. Det fortsatta förfarandet, och särskilt meddelandet av bygglov, grundar sig på denna bedömning. Såsom generaladvokaten anfört i punkt 115 i sitt förslag till avgörande kan den omständigheten att miljökonsekvensbedömningen enligt den slovakiska lagstiftningen görs i ett annat förfarande än det egentliga tillståndsförfarandet, inte medföra en utvidgning av tillämpningsområdet i tiden för direktiv 85/337.
Det framgår även av vad som anförts i punkt 79 i denna dom att stadsplaneringsbeslutet om lokalisering av den deponi som det nationella målet avser utgör en nödvändig förutsättning för att exploatören ska få tillstånd att genomföra det aktuella deponiprojektet. I detta beslut ställs dessutom vissa villkor som exploatören måste uppfylla under genomförandet av projektet.
Domstolen har emellertid, vid prövningen av ett jämförbart förfarande, slagit fast att referensdatumet för fastställande av tillämpningsområdet i tiden för ett direktiv som inför krav på en miljökonsekvensbedömning är det datum då projektet formellt presenterades, eftersom de olika stadierna av projektbedömningen knyter an till varandra så att de utgör ett sammansatt förlopp (dom av den 23 mars 2006, i mål C-209/04, kommissionen mot Österrike, REG 2006, s. I-2755, punkt 58).
Slutligen framgår det av fast rättspraxis att ett tillstånd enligt direktiv 85/337 kan utgöras av en kombination av flera separata beslut när det nationella förfarande som innebär att exploatören får tillstånd att påbörja arbetena för genomförande av sitt projekt består av flera successiva etapper (se, för ett liknande resonemang, dom av den 7 januari 2004 i mål C-201/02, Wells, REG 2004, s. I-723, punkt 52, och av den 4 maj 2006 i mål C-508/03, kommissionen mot Förenade kungariket, REG 2006, s. I-3969, punkt 102). Härav följer att datumet för det formella ingivandet av tillståndsansökan för projektet i så fall är den dag då exploatören gav in en ansökan i syfte att inleda den första etappen av förfarandet.
Mot bakgrund härav kan det konstateras att tillståndsansökan för det deponiprojekt som det nationella målet avser formellt sett ingavs innan det att fristen för införlivande av direktiv 85/337 gick ut. De skyldigheter som följer av detta direktiv är således inte tillämpliga på projektet, varför det saknas anledning att besvara den tredje frågan.
Den fjärde frågan
Den nationella domstolen har ställt den fjärde frågan för att få klarhet i huruvida artiklarna 1 och 15a i direktiv 96/61, i förening med artiklarna 6 och 9 i Århuskonventionen, ska tolkas så, att medlemmarna av den berörda allmänheten, inom ramen för en sådan rättslig prövning som föreskrivs i artikel 15a i direktivet, ska ha rätt att yrka att den domstol eller annat oberoende och opartiskt behörigt organ som inrättats genom lag ska förordna om interimistiska åtgärder i form av inhibition av ett tillstånd enligt artikel 4 i direktivet intill dess att ett slutligt avgörande meddelas.
Medlemsstaterna har, med förbehåll för att de ska iaktta likvärdighetsprincipen och effektivitetsprincipen, i kraft av sin processuella autonomi ett utrymme för skönsmässig bedömning vid genomförandet av artikel 9 i Århuskonventionen och artikel 15a i direktiv 96/61. Det tillkommer dem särskilt att fastställa vilken domstol eller vilket oberoende och opartiskt organ som inrättats genom lag som ska ha behörighet att utföra den rättsliga prövning som avses i dessa bestämmelser, och enligt vilka handläggningsregler denna prövning ska ske, allt under förutsättning att ovannämnda bestämmelser har följts (se, analogt, dom av den 18 oktober 2011 i de förenade målen C-128/09–C-131/09, C-134/09 och C-135/09, Boxus m.fl., REU 2011, s. I-9711, punkt 52).
Det framgår vidare av fast rättspraxis att en domstol som prövar en tvist som ska avgöras utifrån unionsrätten måste kunna bevilja interimistiska åtgärder för att säkerställa den fulla verkan av det senare domstolsavgörandet avseende förekomsten av de rättigheter som gjorts gällande på grundval av unionsrätten (dom av den 19 juni 1990, i mål C-213/89, Factortame m.fl., REG 1990, s. I-2433, punkt 21, svensk specialutgåva, volym 10, s. I-435, och av den 13 mars 2007 i mål C-432/05, Unibet, REG 2007, s. I-2271, punkt 67).
Det ska även tilläggas att rätten att få till stånd en sådan prövning som avses i artikel 15a i direktiv 96/61 ska tolkas mot bakgrund av syftet med detta direktiv. Domstolen har redan slagit fast att detta syfte, såsom det definieras i artikel 1 i direktivet, är att genom samordnade åtgärder förebygga och minska föroreningar som härrör från de verksamheter som anges i bilaga I i luft, vatten och mark, så att en hög skyddsnivå kan uppnås för miljön (dom av den 22 januari 2009 i mål C-437/07, Association nationale pour la protection des eaux et rivières och OABA, REG 2009, s. I-319, punkt 25, och av den 15 december 2011 i mål C-585/10, Møller, REU 2011, s. I-13407, punkt 29).
Nämnda föroreningar skulle emellertid inte kunna förebyggas på ett verkningsfullt sätt genom utnyttjande av rätten att få till stånd en sådan rättslig prövning som avses i artikel 15a i direktiv 96/61 om det vore omöjligt att förhindra fortsatt drift av en anläggning som kan ha beviljats tillstånd i strid med direktivet i avvaktan på ett slutligt avgörande avseende lagenligheten av tillståndet. För att säkerställa att rätten att få till stånd en rättslig prövning enligt artikel 15a i direktivet kan utövas på ett effektivt sätt krävs således att medlemmarna av den berörda allmänheten har rätt att yrka att domstolen, eller det oberoende och opartiska organ som är behörigt, ska förordna om interimistiska åtgärder till förebyggande av dessa föroreningar, såsom i förekommande fall inhibition av det angripna tillståndet
Mot denna bakgrund ska den fjärde frågan besvaras enligt följande: Artikel 15a i direktiv 96/61 ska tolkas så, att medlemmarna av den berörda allmänheten, inom ramen för en sådan rättslig prövning som föreskrivs i denna bestämmelse, ska ha rätt att yrka att den domstol eller annat oberoende och opartiskt behörigt organ som inrättats genom lag ska förordna om interimistiska åtgärder i form av inhibition av ett tillstånd enligt artikel 4 i direktivet intill dess att ett slutligt avgörande meddelas.
Den femte frågan
Den nationella domstolen har ställt den femte frågan för att få klarhet i huruvida ett avgörande från en nationell domstol, som fattats inom ramen för ett nationellt förfarande genom vilket medlemsstaten uppfyller sina åtaganden enligt artikel 15a i direktiv 96/91 och artikel 9.2 och 9.4 i Århuskonventionen och som upphäver ett tillstånd som beviljats i strid med bestämmelserna i nämnda direktiv, kan utgöra ett oberättigat ingrepp i exploatörens äganderätt enligt artikel 17 i Europeiska unionens stadga om de grundläggande rättigheterna.
Mål C‑80/12
Felixstowe Dock and Railway Company Ltd,
Savers Health and Beauty Ltd,
Walton Container Terminal Ltd,
WPCS (UK) Finance Ltd,
AS Watson Card Services (UK) Ltd,
Hutchison Whampoa (Europe) Ltd,
Kruidvat UK Ltd,
Superdrug Stores plc
mot
The Commissioners for Her Majesty’s Revenue and Customs
(begäran om förhandsavgörande från First-Tier Tribunal (Tax Chamber), Förenade kungariket)
Tolkning av artiklarna 43 EG och 48 EG — Etableringsfrihet — Skattelagstiftning — Inkomstskatt för juridiska personer — Skattelättnad — Konsortieyrkande om koncernavdrag (konsortieavdrag) — Nationell lagstiftning som utesluter överföring av underskott inom landet från ett konsortiebolag till ett annat bolag som ingår i en bolagskoncern till vilken ett ’anknytningsbolag’ som också ingår i konsortiet hör — Hemvistkrav för anknytningsbolaget — Diskriminering beroende på platsen för bolagets säte — Yttersta moderbolaget i tredjeland — Kopplingar mellan bolag som löper genom tredjeländer”
I – Inledning
Förenade kungariket tillåter att bolag i skattemässigt hänseende för över underskott till ett annat bolag som det är anknutet till genom vissa kopplingar mellan bolag. Förevarande begäran om förhandsavgörande från First-Tier Tribunal (Tax Chamber) avser i huvudsak frågan huruvida det enligt Europeiska unionens (EU) rättsordning föreligger en inskränkning i etableringsfriheten om sådan överlåtelse av underskott inte får ske när det bolag som utgör anknytningen mellan (i) det bolag som överlåter underskottet och (ii) det bolag som tar över underskottet, har hemvist i en annan medlemsstat. Den hänskjutande domstolen har också frågat huruvida situationen i unionsrättsligt hänseende blir en annan om anknytningen mellan bolag går via bolag i tredjeländer.
Systemet med koncernavdrag i Förenade kungariket medger att underskott överlåts mellan olika bolag i en bolagskoncern ( 2 ) och/eller ett konsortium ( 3 ), vilket därmed möjliggör ett optimalt utnyttjande av dessa underskott i skattehänseende, dock utan att detta leder till att koncernen eller konsortiet konsolideras till en enda ekonomisk enhet i skattehänseende. ( 4 )
Domstolen har än en gång att ta ställning till frågan huruvida den omständigheten att vissa skattskyldiga inte ges tillgång till det i Förenade kungariket gällande systemet för koncernavdrag är förenligt med etableringsfriheten. I målet ICI rörde uteslutandet från systemet med koncernavdrag ett inhemskt holdingbolag som huvudsakligen drev dotterbolag i utlandet, i målet Marks & Spencer avsågs dotterbolag i utlandet och i målet Philips Electronics UK behandlades det i Förenade kungariket belägna fasta driftstället tillhörande ett bolag med hemvist i en annan medlemsstat. ( 5 )
Vad som vid en första anblick skiljer förevarande mål från de tidigare är att kopplingarna mellan bolagen löper via tredjeländer och att det yttersta moderbolaget ( 6 ) har hemvist i ett tredjeland. Denna fråga behöver dock inte vara avgörande för den slutliga bedömningen i förevarande mål av huruvida Förenade kungarikets lagstiftning är förenlig med unionsrätten.
Frågan huruvida unionsrätten aktualiseras i förevarande mål avgörs vidare till viss del av den omständigheten att det i Förenade kungariket är praxis att vederlag utges när underskott överlåts mellan bolag. Detta eftersom förevarande mål grundas på antagandet att ett överlåtande bolag lider en nackdel om det inte kan överlåta underskott till de yrkande bolagen mot vederlag. En sådan ekonomisk nackdel uppkommer endast om det överlåtande bolaget lider en nackdel i fråga om kassaflödet på grund av att det inte kan realisera sitt underskott omedelbart utan att behöva invänta senare räkenskapsår. Om överlåtelsen av underskott sker utan vederlag skulle dock en eventuell nackdel som föranleds av Förenade kungarikets lagstiftning endast märkas på koncernnivå och inte hos det överlåtande bolaget.
II – Nationell rätt, omständigheterna i målet, förfarandet och hänskjutna frågor
A – Förenade kungarikets lagstiftning
De nationella bestämmelser som tillämpats i det nationella målet återfinns i Income and Corporation Taxes Act 1988 (ICTA).
Bolagskoncern” definieras enligt följande i section 413(3) ICTA: Två bolag anses ingå i en koncern om det ena bolaget utgör ett till 75 procent ägt dotterbolag till det andra bolaget eller om båda bolag utgör till 75 procent ägda dotterbolag till ett tredje bolag.
I ICTA föreskrivs två typer av lättnad på koncernnivå: koncernyrkanden avseende koncernavdrag (vilket var i fråga i det ovannämnda målet Marks & Spencer) och konsortieyrkanden avseende koncernavdrag (konsortieavdrag) (vilket var i fråga i de ovannämnda målen ICI och Philips Electronics UK och vilket också är i fråga i förevarande mål).
Enligt section 402 ICTA kan underskott av näringsverksamhet och andra avdragsgilla belopp som får användas för lättnad från inkomstskatt för juridiska personer överlåtas av ett bolag (nedan kallat det överlåtande bolaget) och, på yrkande av ett annat bolag (nedan kallat det yrkande bolaget) medges det yrkande bolaget genom lättnad från inkomstskatt för juridiska personer, så kallat koncernavdrag. I subsection 3 i den bestämmelsen föreskrivs att koncernavdrag, efter framställande av ett så kallat konsortieyrkande, också får medges för bland annat ett överlåtande bolag och ett yrkande bolag när det ena av dem ingår i en koncern och det andra ägs av ett konsortium och ett annat bolag ingår i såväl koncernen som konsortiet.
Enligt subsection 3A i section 402 ICTA medges inte avdrag om inte villkoret i subsection 3B, nämligen att bolaget har hemvist i Förenade kungariket eller saknar hemvist i Förenade kungariket men bedriver verksamhet där via ett fast driftställe, är uppfyllt för såväl det överlåtande som det yrkande bolaget.
I section 406(1) ICTA anges tre definitioner. ”Anknytningsbolag” är ett bolag som ingår i ett konsortium och i en koncern. Ett ”konsortiebolag” är i förhållande till ett anknytningsbolag ett bolag som ägs av det konsortium i vilket anknytningsbolaget ingår. En ”koncernmedlem” är i förhållande till ett anknytningsbolag ett bolag som ingår i den koncern som också anknytningsbolaget ingår i, men som inte själv ingår i det konsortium som anknytningsbolaget ingår i.
I section 406(2) ICTA föreskrivs att ”när anknytningsbolaget … kan framställa ett konsortieyrkande avseende underskott av näringsverksamhet eller ett annat avdragsgillt belopp beträffande ett räkenskapsår för ett bolag som ingår i konsortiet, kan en koncernmedlem framställa ett konsortieyrkande som anknytningsbolaget hade kunnat framställa” motsvarande samma andel av det överlåtna underskottet som om anknytningsbolaget utgjorde det yrkande bolaget.
Det framgår av bestämmelserna i artikel 402(3A) och 402(3B) jämförda med artikel 406(2) ICTA att anknytningsbolaget vad beträffar konsortieyrkanden om koncernavdrag måste ha sitt hemvist i Förenade kungariket eller, om det saknar sådant hemvist, bedriva näringsverksamhet i Förenade kungariket via ett fast driftställe. Anknytningsbolaget ska med andra ord, liksom det överlåtande bolaget och det yrkande bolaget, vara skattskyldiga till inkomstskatt för juridiska personer i Förenade kungariket.
B – Bolagskoncernen och konsortiet
Felixstowe Dock och Railway Company Ltd m.fl. utgör ”de yrkande bolagen”. ( 7 ) De ingår samtliga i Hutchison Whampoa‑koncernen, för vilken det yttersta moderbolaget är Hutchison Whampoa Ltd, ett bolag som bildats i Hongkong där det också har sitt hemvist, och som indirekt äger 100 procent av andelarna i de yrkande bolagen. ( 8 )
Hutchison 3G UK Ltd utgör ”det överlåtande bolaget”. Det ägdes till 100 procent av Hutchison 3G UK Holdings Ltd.
Hutchison 3G UK Holdings Ltd utgjorde konsortiebolaget. Under den relevanta tidsperioden ägdes Hutchison 3G UK Holdings Ltd av ett konsortium bestående av Hutchison 3G UK Investments Sàrl, ett bolag ingående i Hutchison Whampoa‑koncernen som bildats i Luxemburg där det också har sitt hemvist (50,1 procent), tre andra bolag i Hutchison Whampoa‑koncernen som bildats på Brittiska Jungfruöarna där de också har sitt hemvist (totalt 14,9 procent), och två andra bolag som inte har någon anknytning till Hutchison Whampoa‑koncernen (20 procent respektive 15 procent).
Hutchison 3G UK Investments Sàrl utgjorde ”anknytningsbolaget”, och utgjorde länken mellan koncernen och konsortiet. Det var helägt av Hutchison Europe Telecommunications Sàrl, ett bolag som bildats i Luxemburg där det också har sitt hemvist. ( 9 ) Båda bolagen utgör indirekt helägda dotterbolag till Hutchison Whampoa Ltd Ytterligare kopplingar mellan anknytningsbolaget och Hutchison Whampoa Ltd löper genom olika mellanliggande holdingbolag som bildats i Luxemburg och utanför EU/EES (Hongkong, Brittiska Jungfruöarna och Caymanöarna).
C – Det nationella målet och de hänskjutna frågorna
Det överlåtande bolaget bedrev verksamhet som mobiltelefonioperatör. Det ådrog sig betydande kostnader när det installerade sitt system och redovisade därmed stora underskott under de första verksamhetsåren. Vad tillämpningen av section 406(1)(b) ICTA beträffar ägdes det överlåtande bolaget under den aktuella tidsperioden av konsortiebolaget såsom beskrivits ovan.
De yrkande bolagen, vilka redovisade överskott under samma period, önskade utnyttja underskotten i det överlåtande bolaget. Enligt begäran om förhandsavgörande hade det överlåtande bolaget enligt en uppgörelse inom Hutchison Whampoa‑koncernen, rätt till 30 pence för varje 1 GBP av överlåtna underskott. De yrkande bolagen var ”koncernmedlemmar” i den mening som avses i section 406(1)(c) ICTA eftersom de utgjorde indirekta dotterbolag till Hutchison Whampoa Ltd, i vilka sistnämnda bolags andel inte understeg 75 procent. ( 10 )
De yrkande bolagen yrkade konsortieavdrag enligt sections 402(3) och 406 ICTA. Yrkandet avslogs med hänvisning till att anknytningsbolaget (som inte på något sätt var direkt involverat i dessa förfaranden) inte hade hemvist i Förenade kungariket utan i Luxemburg. Det kunde inte överföra någon rätt att yrka konsortieavdrag till något annat bolag i koncernen enligt section 406(1) ICTA eftersom det enligt undantaget i section 402(3B) inte ens för egen del ägde rätt att framställa något sådant yrkande.
Efter det att ärendet överklagats till First-tier Tribunal (Tax Chamber) beslutade denna att vilandeförklara målet och ställa följande frågor till domstolen:
1.
Utgör artiklarna 49 FEUF och 54 FEUF [(tidigare artiklarna 43 EG och 48 EG)] hinder för kravet att anknytningsbolaget ska ha hemvist i Förenade kungariket eller bedriva näringsverksamhet i denna medlemsstat via ett fast driftställe där, när
bestämmelserna i en medlemsstat (såsom Förenade kungariket), innebär att det för att ett bolag (det yrkande bolaget) ska kunna yrka koncernavdrag för underskott i ett bolag som ägs av ett konsortium (konsortiebolag) uppställs som villkor att ett bolag som ingår i samma koncern som det yrkande bolaget också ingår i konsortiet (ett ’anknytningsbolag’), och
moderbolaget i bolagskoncernen (som inte själv utgör det yrkande bolaget, konsortiebolaget eller anknytningsbolaget) inte har sitt säte i Förenade kungariket eller någon annan medlemsstat?
Om den första frågan besvaras jakande: Är Förenade kungariket skyldigt att tillhandahålla ett medel till det yrkande bolaget (till exempel genom att tillåta detta bolag att yrka avdrag för underskott i konsortiebolaget) när
’anknytningsbolaget’ har utövat sin etableringsfrihet men konsortiebolaget och de yrkande bolagen inte har utövat några av de friheter som tillerkänns enligt unionsrätten,
anknytningen mellan det överlåtande bolaget och det yrkande bolaget utgörs av bolag av vilka inte alla är etablerade inom EU/[Europeiska ekonomiska samarbetsområdet (EES)]?”
Skriftliga synpunkter har ingetts av Felixstowe Dock and Railway Company m.fl., den tyska, den franska och den nederländska regeringen samt av Förenade kungarikets regering och Europeiska kommissionen. Förhandling hölls den 3 september 2013, vid vilken samtliga av dessa, med undantag av den franska regeringen, yttrade sig muntligen.
III – Bedömning
A – Inledande anmärkningar
Den hänskjutande domstolens två frågor rör etableringsfriheten. Jag kommer att grunda min bedömning på artiklarna 43 EG och 48 EG, eftersom artiklarna 49 FEUF och 54 FEUF inte är tillämpliga i tiden (ratione temporis) på situationen i det nationella målet.
Jag kommer vid denna bedömning att diskutera de två frågorna tillsammans. Den hänskjutande domstolen har för det första frågat om artiklarna 43 EG och 48 EG, i den situation som är i fråga i det nationella målet, utgör hinder för kravet att anknytningsbolaget, när det gäller systemet med konsortieavdrag, antingen ska ha hemvist i Förenade kungariket eller bedriva näringsverksamhet där via ett fast driftställe. För det andra önskar den hänskjutande domstolen få klarhet i huruvida dessa artiklar innebär ett förbud för en medlemsstat att kräva att det innersta moderbolaget i en bolagskoncern till vilken anknytningsbolaget och de bolag som av skatteskäl tar emot underskotten hör, ska ha hemvist i en medlemsstat eller i en EES-stat, eller att kopplingarna mellan anknytningsbolaget och de bolag som av skatteskäl tar emot underskotten uteslutande utgörs av sådana bolag. Slutligen önskar den hänskjutande domstolen få klarhet i huruvida en sådan åtgärd som den att medge konsortieavdrag för de yrkande bolagen ska finnas att tillgå om Förenade kungarikets bestämmelse utgör ett åsidosättande av etableringsfriheten.
Det ska redan nu klargöras att detta mål inte rör fördelningen av beskattningsrätten mellan medlemsstaterna, även om det enligt vad som framgår av den tyska och den franska regeringens yttranden finns farhågor om att utgången i detta mål kan äventyra deras befogenheter att beskatta internationella bolagskoncerner som kontrolleras av moderbolag med hemvist i tredjeland.
Förevarande mål avser mycket riktigt överlåtelse av underskott från ett bolag som är skattskyldigt till inkomstskatt för juridiska personer i Förenade kungariket, i syfte att kvitta dem mot överskott i ett annat bolag i Förenade kungariket som också är skattskyldigt till inkomstskatt för juridiska personer där. Det är alltså inte fråga om någon gränsöverskridande överlåtelse av underskott mellan bolag med hemvist i olika medlemsstater här, vilket i likhet med vad som var fallet i de ovannämnda målen National Grid Indus ( 11 ) och Philips Electronics UK ( 12 ) skulle aktualisera frågan om fördelningen av beskattningsrätten. Förevarande mål rör endast frågan huruvida det för ett konsortieavdrag får krävas att överlåtelsen av underskott från ett bolag med hemvist i Förenade kungariket till en annan konsortiemedlem får krävas att anknytningsbolaget utgör ett bolag med hemvist i Förenade kungariket eller att det har ett fast driftställe i Förenade kungariket.
I detta sammanhang underlättar det att känna till de tre utvecklingsstadierna beträffande Förenade kungarikets lagstiftning om koncernavdrag. Fram till den 1 april 2000 (det vill säga före den period som är aktuell i förevarande mål), var det inte möjligt att yrka koncernavdrag mellan två systerbolag om deras moderbolag saknade hemvist i Förenade kungariket. Sedan den 1 april 2001 (som är den period som är aktuell i förevarande mål), får bolag som ingår i samma koncern överlåta underskott till varandra oberoende av var moderbolaget har sitt hemvist. Detta innebär att om Hutchison Whampoa‑koncernen (indirekt) hade ägt minst 75 procent av det överlåtande bolaget under den relevanta perioden, i stället för de 65 procent som det faktiskt ägde, så hade det inte förelegat något hinder för de yrkande bolagen att utnyttja det överlåtande bolagets underskott, eftersom sistnämnda bolag ingick i koncernen vid tillämpningen av section 402(1) och 402(2) ICTA. År 2010, efter den period som avses i det nationella målet, har Förenade kungariket ändrat bestämmelserna om koncernavdrag genom Corporation Tax Act 2010, vilket medfört att ett bolag med hemvist i EU/EES kan utgöra anknytningsbolag. Enligt de nya bestämmelserna krävs emellertid att anknytningsbolaget och de yrkande bolagen ingår i samma koncern utan inblandning av ett bolag utanför EU/EES.
Om domstolen följaktligen skulle finna att det föreligger en otillåten restriktion av grundläggande rättigheter kan den nu aktuella lagstiftningen i Förenade kungariket inte motiveras av behovet att upprätthålla fördelningen av beskattningsrätten mellan medlemsstaterna. Inte heller kan behovet av att upprätthålla skattesystemets inre sammanhang åberopas som motivering med hänsyn till den ovan beskrivna utvecklingen av lagstiftningen, som har gjort koncernavdrag möjliga oavsett var moderbolaget eller andra bolag än det överlåtande bolaget och det yrkande bolaget har hemvist. Förenade kungariket har nämligen inte anfört någon motivering för den nationella bestämmelsen i ändrad lydelse eftersom dess ståndpunkt är att det nationella målet inte omfattas av tillämpningsområdet för unionsrätten. ( 13 )
Vidare gäller enligt rättspraxis att även om området för direkt beskattning omfattas av medlemsstaternas behörighet får denna behörighet inte utövas i strid med unionsrätten, närmare bestämt de grundläggande friheter som garanteras i fördragen. Som generaladvokat Kokott har påpekat är medlemsstaterna enligt unionsrätten i princip inte skyldiga att i sina respektive lagstiftningar om inkomstskatt för juridiska personer föreskriva en rätt till koncernavdrag för underskott. Utformningen av skattesystemet ankommer nämligen på medlemsstaterna själva. I den mån en sådan rättighet medges ska den emellertid tillämpas på ett sätt som är förenligt med de grundläggande friheterna enligt unionsrätten, i synnerhet etableringsfriheten. ( 14 )
B – Det sätt på vilket koncernavdraget fungerar
I ekonomiska termer möjliggör det slags koncernavdrag som är tillämpligt i Förenade kungariket för det överlåtande bolaget att föra över sina underskott till det yrkande bolaget, som kan dra av dem från sitt skattepliktiga överskott. Detta medför att det överlåtande bolaget förlorar rätten att utnyttja dessa underskott vid beskattningen, närmare bestämt möjligheten att spara underskotten till kommande räkenskapsår. ( 15 )
Praxis i Förenade kungariket synes vara att denna överlåtelse sker mot vederlag, ( 16 ) vilket ofta motsvarar värdet av den inkomstskatt för juridiska personer som sparas in tack vare underskottet, även om detta vederlag saknar stöd i lagstiftningen, eventuellt med förbehåll för det fallet att de bolagsrättsliga förvaltningsskyldigheter som åvilar det överlåtande bolagets ledning för med sig ett sådant krav. Exempelvis har de yrkande bolagen i förevarande fall gått med på att betala 30 pence per 1 GBP för överlåtna underskott.
Eftersom Förenade kungarikets system med koncernavdrag inte baseras på skattemässig konsolidering på koncernnivå av över- och underskott, står det klart att ett överlåtande bolag i egenskap av självständig juridisk person med vinstsyfte normalt sett inte skulle gå med på att utan vederlag överlåta underskott som det senare skulle kunna använda för att minimera sina egna framtida skatter. Genom att överlåta underskotten mot vederlag som återspeglar den tillämpliga inkomstskattesatsen för juridiska personer, monetäriserar det överlåtande bolaget sina underskott på ett tidigare (och säkrare) stadium, vilket leder till en kassaflödesfördel.
Om existerande praxis i Förenade kungariket skulle vara en annan än den ovan beskrivna, vore det svårt att se varför ett överlåtande bolag skulle lida någon egentlig skada på grund av en bestämmelse i lag som hindrar det från att överlåta sina underskott till ett annat bolag, det vill säga från att överlåta tillgångar som kan ha ett ekonomiskt värde i form av underlag för kvittning vid framtida beskattning till en utomstående mot ett vederlag som inte återspeglar deras värde för det överlåtande bolaget. Det skulle också vara svårt att hävda att en bestämmelse i lag som hindrar ett bolag med vinstsyfte från att överlåta sina tillgångar utan vederbörligt vederlag skulle utgöra en inskränkning av etableringsfriheten. Utan dessa faktiska omständigheter skulle därmed de nackdelar som följer av lagstiftningen i Förenade kungariket inte märkas för det överlåtande bolaget utan endast för de bolag som befinner sig högre upp i koncernen och konsortiet än det överlåtande bolaget och de yrkande bolagen, det vill säga på koncernnivå i form av en högre skattebörda för koncernen som helhet.
Denna kassaflödesfördel, eller möjligheten att vinna en sådan fördel, bör öka värdet på det överlåtande bolaget och därmed även på andelsinnehav i bolaget. Detta innebär att möjligheten till koncernavdrag gynnar ägarna i det överlåtande bolaget, oavsett om dessa utgör direkta eller indirekta moderbolag, eller konsortiemedlemmar med minoritetsägande. ( 17 )
För ett yrkande bolag är en sådan lösning ekonomiskt neutral: det betalar ett belopp till det överlåtande bolaget som motsvarar den skatt det undviker tack vare överlåtelsen i stället för att betala samma belopp till skatteförvaltningen. Eftersom det emellertid enligt Förenade kungarikets lagstiftning krävs att det yrkande bolaget och anknytningsbolaget tillhör samma koncern, vilket även gäller i fråga om konsortieavdrag, förklaras arrangemangen mellan de yrkande bolagen och de överlåtande bolagen av den fördel som koncernen vinner genom koncernavdraget, eftersom det leder till en lägre skattebörda på koncernnivå. ( 18 )
C – Vilken grundläggande frihet är relevant i materiellt hänseende?
När det gäller de kriterier som slagits fast i domstolens praxis kan det framstå som tveksamt huruvida Förenade kungarikets lagstiftning har att göra med etableringsfriheten. Etableringsfrihetens tillämplighet avgörs enligt domstolen av graden av kontroll som utövas över ett visst bolag. I förevarande mål kan graden av kontroll som krävs enligt nationell rätt vara allt från 5 procent, vilket knappast ger ”kontroll”, till 74,99 procent. Svaret på denna fråga tycks emellertid framgå av omständigheterna i målet vilket jag ämnar förklara nedan, och det är också etableringsfriheten som den hänskjutande domstolen har hänvisat till när den ställt sina frågor.
Tredjelandsaspekter som har att göra med den komplicerade bolagsstrukturen i Hutchison Whampoa‑koncernen ger upphov till frågan huruvida den relevanta lagstiftningen i Förenade kungariket ska bedömas mot bakgrund av etableringsfriheten, som inte är tillämplig i förhållande till tredjeländer, och/eller mot bakgrund av den fria rörligheten för kapital, som är tillämplig även i förhållande till tredjeländer.
Domstolen slog i sin dom av den 13 november 2012 i mål C‑35/11, Test Claimants in the FII Group Litigation, fast att frågan huruvida en nationell lagstiftning omfattas av den ena eller andra fria rörligheten enligt numera fast rättspraxis ska avgöras med beaktande av ändamålet med den aktuella lagstiftningen. En nationell lagstiftning som endast ska tillämpas på andelsinnehav som ger ett bestämmande inflytande över ett bolags beslut och verksamhet, omfattas etableringsfriheten. Däremot ska de nationella bestämmelser som är tillämpliga på andelsinnehav som förvärvats uteslutande i placeringssyfte utan avsikt att erhålla något inflytande på förvaltning och kontroll av företaget bedömas enbart utifrån den fria rörligheten för kapital. ( 19 )
I situationer där det inte är möjligt att utifrån ändamålet med den nationella lagstiftningen fastställa huruvida denna till övervägande del omfattas av artikel 49 FEUF eller artikel 63 FEUF, tar domstolen hänsyn till faktiska omständigheter i det enskilda fallet i syfte att avgöra om den situation som tvisten i det nationella målet avser omfattas av den ena eller andra av dessa bestämmelser (min kursivering). ( 20 )
Här ska en distinktion göras mellan de två typerna av koncernavdrag som Förenade kungarikets lagstiftning erbjuder. Ur ett ändamålsperspektiv tar Förenade kungarikets bestämmelser om koncernyrkande om koncernavdrag klart sikte på de andelsinnehav som ger aktieägaren ett bestämmande inflytande över ett bolags beslut och verksamhet. De är tillämpliga på bolag som till minst 75 procent utgör dotterbolag. Bestämmelserna omfattas därmed av etableringsfriheten.
När det gäller konsortieyrkanden om koncernavdrag är situationen mera oklar. Bestämmelser om konsortieavdrag är tillämpliga i situationer där minst 75 procent av kapitalet i konsortiebolaget ägs av konsortiemedlemmar, vilka var för sig inte får äga mindre än 5 procent och inte 75 procent eller mer. ( 21 ) Detta omfattar situationer där det finns en dominerande ägare men också situationer där det finns många sinsemellan fristående aktieägare. I teorin skulle det kunna finnas ett konsortiebolag med 20 andelsägare som var och en äger 5 procent i konsortiebolaget. Detta skulle kunna ge upphov till en situation med 20 anknytningsbolag där konsortiebolaget skulle kunna överlåta sina underskott, i femprocentiga delar, till 20 olika bolagskoncerner.
Enligt min mening är Förenade kungarikets bestämmelser om konsortieavdrag inte avsedda att enbart tillämpas på de andelsinnehav som ger innehavaren rätt att utöva ett bestämmande inflytande över ett bolags beslut. Som ombudet för de yrkande bolagen anförde under förhandlingen, innehåller inte Förenade kungarikets lagstiftning något krav på att konsortiemedlemmarna utövar någon slags legaldefinierad kollektiv kontroll över konsortiebolaget. ( 22 ) Holdingbolag som får beaktas vid konsortieavdrag kan därför enligt min mening betraktas som direkta investeringar och eventuella inskränkningar för dem kan anses utgöra restriktioner för fria kapitalrörelser. ( 23 )
Förenade kungarikets bestämmelser tillåter emellertid även situationer där konsortiebolaget kontrolleras av en enda bolagskoncern. Detta är fallet beträffande det överlåtande bolaget i förevarande mål: 65 procent av det bolaget ägs indirekt av Hutchison Whampoa‑koncernen (50,1 procent via anknytningsbolaget och 14,9 procent via tre koncernbolag på Brittiska Jungfruöarna). De aktuella bestämmelserna kan följaktligen innebära en inskränkning i etableringsfriheten och den situation som är i fråga i det nationella målet bör anses ingå i tillämpningsområdet för denna grundläggande frihet.
Jag anser mot bakgrund av dessa överväganden att omständigheterna i målet faller inom tillämpningsområdet för artikel 43 EG, vilket innebär att Förenade kungarikets system med koncernavdrag i första hand ska prövas mot etableringsfriheten.
D – Huruvida det föreligger en inskränkning av etableringsfriheten
Den etableringsfrihet som enligt artikel 43 EG tillerkänns unionsmedborgare, och som för dem innefattar en rätt att starta och utöva verksamhet som egenföretagare samt rätt att bilda och driva företag på de villkor som etableringslandets lagstiftning föreskriver för egna medborgare, inbegriper i enlighet med artikel 48 EG en rätt för bolag som bildats i överensstämmelse med en medlemsstats lagstiftning, och som har sitt säte, sitt huvudkontor eller sin huvudsakliga verksamhet inom Europeiska unionen, att utöva verksamhet i den berörda medlemsstaten genom ett dotterbolag, en filial eller ett kontor. Då det uttryckligen anges i artikel 43 första stycket andra meningen EG att ekonomiska aktörer fritt ska kunna välja den juridiska form som är lämplig för att bedriva verksamhet i en annan medlemsstat, får detta fria val inte begränsas i den mottagande medlemsstaten genom diskriminerande skattebestämmelser. ( 24 )
Enligt Förenade kungarikets lagstiftning ska anknytningsbolaget ha hemvist i Förenade kungariket eller, om det saknar hemvist där, bedriva verksamhet i den medlemsstaten via ett fast driftställe. Denna bestämmelse utgör en klar inskränkning av etableringsfriheten för anknytningsbolaget, som har hemvist i Luxemburg, och dess direkta moderbolag, som också har hemvist i Luxemburg.
Domstolen fann i sin dom i det ovannämnda målet Marks & Spencer att ”[e]tt sådant koncernavdrag som är i fråga i målet vid den nationella domstolen innebär en skattelättnad för de berörda bolagen. Koncernavdraget innebär ett tidigare utnyttjande av förluster i bolag som dras med underskott genom att förlusterna omedelbart kan utnyttjas mot vinster i andra koncernbolag och medför således en [likviditetsfördel] för koncernen.” ( 25 ) Innebär detta att nackdelen upplevs endast på koncernnivå, eller av det yttersta moderbolaget, som i förevarande fall är ett företag i tredjeland? Jag anser inte att så är fallet.
Som jag har förklarat ovan innebär Förenade kungarikets system med koncernavdrag i faktiskt hänseende att över- och underskott kvittas inom en koncern och/eller ett konsortium, inte genom en konsoliderad skattemässig redovisning eller genom en överföring av skattepliktigt överskott i form av ett koncernbidrag, utan som en ordning där underskott överlåts mot vederlag, vilket innebär en kassaflödesfördel för det överlåtande bolaget. Om överlåtelse av underskott inte tillåts, och därmed inte heller konsortieavdrag, på grund av anknytningsbolagets hemvist, är det i första hand det överlåtande bolaget som lider en ekonomisk nackdel genom att det går miste om en kassaflödesfördel. I domstolens praxis har en sådan kassaflödesnackdel ansetts utgöra en oförmånlig behandling som kan utgöra en inskränkning. ( 26 ) Nackdelar som ett bolag lider på grund av moderbolagets hemvist ansågs i domen i de förenade målen Metallgesellschaft m.fl. vara tillräckligt för att utgöra ett åsidosättande av etableringsfriheten. ( 27 )
Denna nackdel är också märkbar för ägarna till det överlåtande bolaget i form av ett lägre värde på deras andelsinnehav, oberoende av om dessa utgör kontrollinnehav, stabila minoritetsinvesteringar eller portföljinvesteringar. Det är naturligtvis endast den förstnämnda kategorin som är relevant när det gäller etableringsfriheten.
I förevarande mål förfördelas alltså anknytningsbolaget med hemvist i Luxemburg, vilket indirekt äger 50,1 procent av det överlåtande bolaget med hemvist i Förenade kungariket, mindre i förhållande till ett bolag med hemvist i Förenade kungariket, vilket befinner sig i en jämförbar situation, när det gäller dess förmåga att utgöra anknytning mellan de två bolagen i Förenade kungariket, vilka är skattskyldiga till inkomstskatt för juridiska personer där. Den omständigheten att nackdelen också återspeglas i värdet på det luxemburgska anknytningsbolaget och därför även är märkbart för dess ägare, vilka delvis utgörs av bolag med hemvist i tredjeland, och i slutändan av det yttersta moderbolag som kontrollerar den komplicerade bolagsstrukturen, ändrar inte detta.
Det är därför fråga om direkt diskriminering på grund av anknytningsbolagets nationalitet. Förenade kungarikets bestämmelser leder till att det är förmånligare för anknytningsbolagets moderbolag att placera sitt dotterbolag i Förenade kungariket än i något annat land.
Som jag har förklarat ovan har inte Förenade kungarikets regering anfört några grunder som kan motivera den inskränkning som den nationella lagstiftningen medför. Jag kan därför inte ta ställning till den frågan här.
I detta skede bör det också utrönas huruvida de yrkande bolagen faktiskt har rätt att åberopa etableringsfriheten. Det framgår klart av domen i det ovannämnda målet Philips Electronics UK ( 28 ) att bolag i skattehänseende kan åberopa inskränkningar i etableringsfriheten för ett annat bolag som är anknutet till förstnämnda bolag i den mån dessa inskränkningar påverkar deras egen beskattning. Den omständigheten att varken det överlåtande bolaget eller de yrkande bolagen själva har utövat sin etableringsfrihet är således irrelevant i detta avseende.
De yrkande bolagen kan därför för sin egen beskattning åberopa den inskränkning för etableringsfriheten som gäller för anknytningsbolaget i den mån Förenade kungarikets bestämmelser, sådana de tolkas av den nationella domstolen, är oförenliga med artiklarna 43 EG och 48 EG.
Min slutsats så långt är att kravet på att anknytningsbolaget ska ha hemvist eller ett fast driftställe i Förenade kungariket för att ett konsortieyrkande om koncernavdrag ska vara möjligt utgör en inskränkning av etableringsfriheten som inte kan motiveras och att kravet därför är otillåtet enligt artiklarna 43 EG och 48 EG.
E – Tredjeländer och etableringsfriheten
Etableringsfrihetens förhållande till tredjeländer är viktigt i förevarande fall eftersom den hänskjutande domstolen med sin andra fråga önskar få klarhet i huruvida Förenade kungariket är skyldigt att erbjuda medel för det yrkande bolaget genom att exempelvis låta det bolaget yrka avdrag för underskott i konsortiebolaget, när anknytningsbolaget har utövat sin etableringsfrihet men konsortiebolaget och de bolag som framställt yrkandena inte har utövat någon av de friheter som hägnas av unionsrätten, och anknytningen mellan det överlåtande bolaget och det yrkande bolaget utgörs av bolag av vilka inte samtliga har hemvist i EU/EES.
Denna fråga ska enligt min mening bedömas mot bakgrund av den första frågan eftersom den i allt väsentligt avser det materiella innehållet i etableringsfriheten, och inte de medel som står till buds i processuell mening enligt denna frihet. ( 29 ) Skulle det med andra ord fortfarande vara tillåtet att kräva att anknytningsbolaget är ett bolag i EU/EES eller att kedjan mellan det överlåtande bolaget och de yrkande bolagen inte inbegriper bolag i tredjeland, även när fördraget innebär ett hinder för kravet att anknytningsbolaget antingen ska ha hemvist i Förenade kungariket eller ett fast driftställe där?
Till skillnad från den fria rörligheten för kapital är etableringsfriheten inte tillämplig i förhållande till tredjeländer. Innebär detta att bolag i EU som i själva verket kontrolleras av bolag i tredjeländer eller av fysiska personer inte omfattas av etableringsfriheten? Påverkas med andra ord det luxemburgska anknytningsbolagets etableringsfrihet av att det kontrolleras av ett moderbolag i tredjeland?
Det ska här erinras om att artikel 48 EG likställer bolag som bildats i överensstämmelse med en medlemsstats lagstiftning och som har sitt säte, sitt huvudkontor eller sin huvudsakliga verksamhet inom Europeiska unionen med fysiska personer som är medborgare i medlemsstaten såvitt gäller etableringsfriheten. Som domstolen slog fast i sin dom i det ovannämnda målet ICI ( 30 ) är det bolagets säte i den mening som avses i artikel 48 EG som knyter bolaget till rättssystemet i en viss stat, på samma sätt som medborgarskapet för juridiska personer.
Det finns inte något stöd i fördraget eller i domstolens praxis för att den etableringsfrihet som bolagen i artikel 48 EG åtnjuter enligt unionsrätten skulle begränsas eller påverkas för de bolag som kontrolleras av juridiska eller fysiska personer i ett tredjeland. Bedömningen att ett bolag har hemvist i unionen baseras på var sätet är beläget och på den rättsordning enligt vilken bolaget har bildats, och inte på var aktieägarna har hemvist eller är medborgare. Om bolag med hemvist i unionen inte skulle omfattas av denna frihet, skulle många juridiska personer vars säte är beläget i Europeiska unionen utestängas från etableringsfriheten, och medlemsstater skulle även i annat fall, och då inte bara vid beskattningen, kunna diskriminera dem.
Domen i målet Halliburton Services ( 31 ) visade att de rättigheter som bolagen i medlemsstaterna åtnjuter enligt unionsrätten inte påverkades av att deras moderbolag, Halliburton Inc., hade hemvist i Amerikas förenta stater. Några längre gående slutsatser kan dock inte dras av denna dom när det gäller situationer där bolag i unionen utan gemensamt moderbolag i unionen ingår i en bolagskoncern utanför unionen. I domen i det ovannämnda målet Halliburton Services hade den nationella domstolen redan slagit fast att enligt det bilaterala skatteavtalet mellan Nederländerna och Amerikas förenta stater fick inte det nederländska dotterbolag som köpt det tyska dotterbolagets nederländska fasta driftställe diskrimineras på grund av att koncernens moderbolag bildats i Förenta staterna. ( 32 )
I förevarande fall åtnjuter därför det i Luxemburg registrerade anknytningsbolaget och dess direkta moderbolag, som också är registrerat i Luxemburg, etableringsfrihet och detta oberoende av att de ytterst kontrolleras av ett moderbolag med hemvist i Hongkong.
F – Tillåtna inskränkningar
Innebär detta att Förenade kungariket inte får kräva att det ska finnas en obruten kedja inom EU/EES mellan det överlåtande bolaget och de yrkande bolagen? Kommissionen har i sina yttranden hävdat att Förenade kungariket skulle tillämpa ett sådant krav men att så inte skedde under den period som är aktuell i det nationella målet.
Jag anser inte att den situationen leder till att denna aspekt av den hänskjutande domstolens frågor blir hypotetiska eller medför att frågan om tredjeländer blir irrelevant på så sätt att den inte ska beaktas av domstolen. I en situation där en nationell bestämmelse innebär en diskriminering av ”utländska” juridiska eller fysiska personer, varför den är att anse som oförenlig med unionsrätten, är det nämligen inte otänkbart att en nationell domstol skulle kunna åtgärda den situationen genom en tolkning som innebär att sådan diskriminering av medborgare eller bolag i EU/EES undanröjs utan att fördelen i form av integrering utsträcks till juridiska eller fysiska personer i tredjeland. Huruvida detta är rättsligt möjligt får avgöras enligt nationell rätt. Unionsrätten innehåller inte något krav på att andra grundläggande friheter än fri rörlighet för kapital utsträcks till subjekt i tredjeland. ( 33 )
I domen i målet Test Claimants in the Thin Cap Group Litigation ( 34 ) slog domstolen fast att situationer där moderbolaget, som kontrollerar långivande och låntagande bolag, har hemvist i en stat som inte utgör en medlemsstat, inte omfattas av etableringsfriheten. Domstolen fann att behandlingen av ränta som det låntagande bolaget betalade som utdelning inverkade på etableringsfriheten, men endast beträffande moderbolaget i tredjeland som hade en viss kontroll över vart och ett av bolagen, vilket gav det möjlighet att påverka valet av finansieringsform för dessa bolag. I en sådan situation var artiklarna 43 EG och 48 EG inte tillämpliga.
Eftersom etableringsfriheten inte sträcker sig till tredjeländer hindrar inte unionsrätten att Förenade kungariket uppställer ett krav i sin lagstiftning på att anknytningsbolaget ska vara etablerat i EU/EES. Om alltså det överlåtande bolaget, när det gäller konsortieavdrag, inte får överlåta underskott när det berörda anknytningsbolaget är ett bolag i tredjeland, omfattas alltså inte situationen av tillämpningsområdet för artikel 43 EG. Om exempelvis anknytningsbolaget i det nationella målet, som både ingår i konsortiet och i koncernen, hade bildats på Brittiska Jungfruöarna i stället för i Luxemburg, skulle dess etableringsfrihet inte kunna åberopas till stöd för ett yrkande om konsortieavdrag. Detta skulle vara fallet även om moderbolaget till bolaget med hemvist på Brittiska Jungfruöarna i sin tur har hemvist i EU/EES.
Jag har ovan förordat en tolkning som å ena sidan innebär att etableringsfriheten åsidosätts när möjligheten att överlåta underskott utesluts på grund av att anknytningsbolaget är ett bolag i EU/EES men å andra sidan att det inte är fråga om något åsidosättande när anknytningsbolaget är ett bolag i tredjeland. Vid denna tolkning har jag prövat konsortieavdragssystemet ur det överlåtande bolagets perspektiv och de nackdelar det kan lida, vilket när det gäller etableringsfriheten påverkar bolagets ägare. Problemet måste också belysas ur de yrkande bolagens perspektiv.
Enligt Förenade kungarikets lagstiftning krävs att de yrkande bolagen tillhör samma koncern som anknytningsbolaget, vilket innebär att det yrkande bolaget måste utgöra ett till 75 procent ägt dotterbolag till anknytningsbolaget eller vice versa, eller så måste båda bolagen utgöra till 75 procent ägda dotterbolag till ett tredje bolag. I förevarande fall utgör anknytningsbolaget och de yrkande bolagen helägda dotterbolag till Hutchison International Limited, ett bolag i Hongkong som i sin tur utgör ett helägt dotterbolag till det yttersta moderbolaget i koncernen, Hutchison Whampoa Ltd Kedjorna från anknytningsbolaget och de yrkande bolagen till deras gemensamma moderbolag går via bolag i EU/EES såväl som via bolag i tredjeländer. De har inte något gemensamt moderbolag i EU/EES.
I ett sådant system som det i Förenade kungariket gällande konsortieavdraget, kan nationella bestämmelser om den erforderliga länken mellan anknytningsbolaget och det yrkande bolaget påverka etableringsfriheten för deras innersta gemensamma moderbolag, vilket åtnjuter den ekonomiska fördel som skapas genom möjligheten att kvitta underskott i ett bolag mot ett skattepliktigt överskott i ett annat bolag, vilket minskar det sammanlagda beskattningsunderlaget för dess (under)koncern. Om det innersta gemensamma moderbolaget är ett bolag i EU/EES, kan nationella anknytningsbestämmelser skapa otillåtna inskränkningar av etableringsfriheten. Om detta innersta gemensamma moderbolag är ett företag i tredjeland, faller situationen utanför tillämpningsområdet för etableringsfriheten vilket följer av domen i det ovannämnda målet Test Claimants in the Thin Cap Group Litigation.
Vidare gäller att om kedjan mellan det innersta gemensamma moderbolaget i EU/EES och anknytningsbolaget respektive de yrkande bolagen löper via tredjeländer, faller situationen utanför tillämpningsområdet för artiklarna 43 EG och 48 EG. Etableringsfriheten utsträcker inte rätten att bilda dotterbolag eller filialer i medlemsstater till juridiska personer i tredjeländer. Liksom nationaliteten för aktieägare med kontrollinnehav saknar betydelse för huruvida bolag i EU/EES åtnjuter etableringsfrihet, saknar den också betydelse för frågan om denna frihet inte föreligger för bolag i tredjeländer.
G – Fri rörlighet för kapital
Som jag har förklarat ovan är det möjligt att de relevanta bestämmelserna i Förenade kungariket om konsortielättnad kan eller bör anses påverka den fria rörligheten för kapital, närmare bestämt direkta investeringar i anknytningsbolagets kapital. Jag anser inte att detta ändrar utgången av min ovan redovisade bedömning såvitt avser förhållanden inom EU/EES. Hindret mot att överlåta underskott skapar nämligen även nackdelar för dem som äger andelar i anknytningsbolaget oberoende av om de innehar kontrollposter eller mindre poster.
Om den fria rörligheten för kapital påverkas kommer detta att kräva att tillämpningsområdet för Förenade kungarikets koncernavdrag utsträcks till att även gälla för bolag i tredjeländer. Eftersom Förenade kungarikets lagstiftning även uteslöt anknytningsbolag i tredjeländer från tillämpningsområdet för konsortieavdrag före den 31 december 1993, skulle de relevanta bestämmelserna till följd av standstill-klausulen i artikel 57.1 EG (nu artikel 64.1 FEUF) inte träffas av förbudet mot restriktioner för fria kapitalrörelser. ( 35 )
H – Förslag till svar
Jag föreslår därför att den första frågan besvaras enligt följande. Under sådana förhållanden som de i målet vid den hänskjutande domstolen aktuella, utgör artiklarna 43 EG och 48 EG hinder för ett krav som när det gäller systemet med konsortieavdrag innebär att anknytningsbolaget antingen ska ha hemvist i den berörda medlemsstaten eller bedriva näringsverksamhet i den medlemsstaten via ett där beläget fast driftställe. Dessa artiklar utgör emellertid inte hinder för en medlemsstat att kräva att det innersta gemensamma moderbolaget i den bolagskoncern som anknytningsbolaget och de bolag som för skatteändamål övertar underskotten tillhör, ska vara ett bolag i EU/EES och att kopplingar mellan anknytningsbolaget och de bolag som för skatteändamål övertar underskotten uteslutande utgörs av bolag i EU/EES. Vad gäller den andra frågan räcker det att besvara denna på samma sätt som den fjärde frågan i det ovannämnda målet Philips Electronics UK.
IV – Förslag till avgörande
Mot bakgrund av ovan redovisade överväganden föreslår jag att domstolen ska besvara frågorna från First-Tier Tribunal (Tax Chamber) enligt följande.
Under sådana förhållanden som de i målet vid den hänskjutande domstolen aktuella, utgör artiklarna 43 EG och 48 EG (nu artiklarna 49 FEUF och 54 FEUF) hinder för ett krav som när det gäller systemet med konsortieavdrag innebär att anknytningsbolaget antingen ska ha hemvist i den berörda medlemsstaten eller bedriva näringsverksamhet i den medlemsstaten via ett där beläget fast driftställe. Dessa artiklar utgör emellertid inte hinder för att i nationell lagstiftning kräva att det innersta gemensamma moderbolaget i den bolagskoncern som anknytningsbolaget och de bolag som för skatteändamål övertar underskotten tillhör, ska ha hemvist i en av medlemsstaterna eller i ett land som tillhör Europeiska ekonomiska samarbetsområdet, och att kopplingar mellan anknytningsbolaget och de bolag som för skatteändamål övertar underskotten uteslutande utgörs av sådana bolag.
Den nationella domstolen ska underlåta att tillämpa varje bestämmelse i den nationella lagstiftningen som strider mot artiklarna 43 EG och 48 EG.
Originalspråk: engelska.
I det här aktuella sammanhanget avses med bolagskoncern moderbolag och dotterbolag i form av en ekonomisk enhet som står under gemensam kontroll.
Ett konsortium kan generellt karaktäriseras som en sammanslutning av två eller flera bolag i syfte att delta i en gemensam verksamhet eller att gemensamt dela resurser för att uppnå ett gemensamt mål. Enligt skattelagstiftningen i Förenade kungariket krävs emellertid för ett konsortium att ett visst minsta ägande ska uppnås, dock utan krav på något gemensamt mål.
Se generaladvokaten Poiares Maduros förslag till avgörande i mål C-446/03, Marks & Spencer (REG 2005, s. I-10837), punkt 17.
Dom av den 16 juli 1998 i mål C-264/96, ICI (REG 1998, s. I-4695), av den 13 december 2005 i mål C-446/03, Marks & Spencer (REG 2005, s. I-10837), och av den 6 september 2012 i mål C‑18/11, Philips Electronics UK.
I förevarande mål ska det skiljas mellan begreppen ”innersta gemensamma moder(bolag)” och ”yttersta moder(bolag)”. Det förra kan beskrivas på följande sätt: Bolag C är det innersta gemensamma moderbolaget i förhållande till bolagen A och B om A och B utgör dess direkta eller indirekta dotterbolag och bolag C inte har något dotterbolag D som skulle utgöra moderbolag till såväl bolag A som bolag B. Det yttersta moderbolaget i en bolagskoncern är ett bolag som utgör direkt eller indirekt moderbolag för samtliga koncernbolag men som inte självt utgör dotterbolag till något annat bolag.
De yrkande bolagen är: Felixstowe Dock and Railway Company Ltd, Savers Health and Beauty Ltd, Walton Container Terminal Ltd, WPCS (UK) Finance Ltd, AS Watson Card Services (UK) Ltd, Hutchison Whampoa (Europe) Ltd, Kruidvat UK Ltd och Superdrug Stores plc.
Relevanta subjekt mellan Hutchison Whampoa Ltd och de yrkande bolagen utgjordes av olika mellanliggande holdingbolag som bildats utanför EU/EES (Hongkong eller Brittiska Jungfruöarna) och i EU (Förenade kungariket eller Nederländerna).
Ett bolag i Hutchison Whampoa‑koncernen förvärvade sedermera (den 23 juni 2005) de två sistnämnda bolagen, varigenom också 3G UK holdings Ltd kom att ingå i koncernen enligt definitionen i section 413(3)(a) ICTA.
Enligt section 413(3) ICTA.
Dom av den 29 november 2011 i mål C‑371/10, National Grid Indus (REU 2011, s. I-12273), punkt 45.
Punkt 23. Andra mål där frågan om fördelningen av beskattningsrätten uppkommit är till exempel det ovannämnda målet Marks & Spencer, domen, punkt 45, dom av den 15 maj 2008 i mål C-414/06, Lidl Belgium (REG 2008, s. I-3601), punkt 31, av den 25 februari 2010 i mål C‑337/08, X Holding (REU 2010, s. I‑1215), punkt 28, och av den 21 februari 2013 i mål C‑123/11, A Oy, punkt 23.
Den nederländska regeringen anser däremot att det föreligger en inskränkning av etableringsfriheten som kan motiveras.
Se generaladvokaten Kokotts förslag till avgörande i det ovannämnda målet Philips Electronics UK, punkt 22 och där angiven rättspraxis.
Se generaladvokaten Poiares Maduros förslag till avgörande i det ovannämnda målet Marks & Spencer, punkt 15.
Se generaladvokaten Kokotts förslag till avgörande i det ovannämnda målet Philips Electronics UK, punkterna 14 och 29.
Att en kassaflödesnackdel på koncernnivå kan innebära en inskränkning av etableringsfriheten underströks av generaladvokaten Sharpston i hennes förslag till avgörande i det ovannämnda målet Lidl Belgium, punkterna 29 och 30.
Domstolen erkände denna fördel på koncernnivå i domen i det ovannämnda målet Marks & Spencer, punkt 32 (se nedan för citat).
Dom av den 13 november 2012 i mål C‑35/11, Test Claimants in the FII Group Litigation, punkterna 90–92.
Domen i det ovannämnda målet Test Claimants in the FII Group Litigation, punkterna 93 och 94.
Se sections 402(3), 406(1) och 413(6) ICTA.
Detta till skillnad från domen av den 24 maj 2007 i mål C-157/05, Holböck (REG 2007, s. I-4051), där det var fråga om gemensam kontroll över ett bolag av andelsägare utan kontroll.
Det ska här erinras om att investeringar som ger kontroll alltid utgör direkta investeringar, men att det också finns investeringar som inte ger kontroll men som inte heller är rent ekonomiska, det vill säga portföljinvesteringar, eftersom dessa är avsedda att åstadkomma stabila förhållanden vad gäller målbolaget. När det gäller direkta investeringar enligt unionsrätten, har domstolen slagit fast att artikel 63 FEUF om fri rörlighet för kapital i princip omfattar kapitalrörelser som innebär en etablering eller direkta investeringar. Sistnämnda begrepp avser en form av andelsinnehav i ett företag genom innehav av aktier som ger möjlighet att faktiskt ta del i kontrollen och ledningen av företaget (se dom av den 17 september 2009 i mål C-182/08, Glaxo Wellcome (REG 2009, s. I-8591), punkt 40, av den 21 oktober 2010 i mål C‑81/09, Idrima Tipou (REU 2010, s. I‑10161), punkt 48, och domen i det ovannämnda målet Test Claimants in the FII Group Litigation, punkt 102). I OECD‑termer avser direkta investeringar ändamålet att åstadkomma ett bestående ägande. Detta betyder bland annat att det ska föreligga ett långsiktigt förhållande och en betydande grad av inflytande över ledningen av företaget. Det direkta eller indirekta ägandet om 10 procent eller mer av rösterna påvisar ett sådant förhållande. Se OECD Benchmark Definition of Foreign Direct Investment, fjärde utgåvan 2008, s. 48, punkt 117, och Modell för skatteavtal beträffande inkomst och förmögenhet, förkortad version 2010 (tillgänglig på engelska på www.oecd.org). Se även Smit, D., EU Freedoms, Non-EU Countries and Company Taxation, Kluwer Law International, 2012, sidorna 64 och 68.
Domen i det ovannämnda målet Philips Electronics UK, punkterna 12 och 13.
Domen i det ovannämnda målet Marks & Spencer, punkt 32.
Dom av den 12 december 2006 i mål C-446/04, Test Claimants in the FII Group Litigation (REG 2006, s. I-11753), punkt 84.
Dom av den 8 mars 2001 i de förenade målen C-397/98 och C-410/98, Metallgesellschaft m.fl. (REG 2001, s. I-1727), punkt 43.
Punkt 39.
Se generaladvokaten Kokotts förslag till avgörande i det ovannämnda målet Philips Electronics UK, punkt 81.
Punkt 20.
Dom av den 12 april 1994 i mål C-1/93, Halliburton Services (REG 1994, s. I-1137; svensk specialutgåva, volym 15, s. 71).
Se punkt 6 i domen.
Situationen här skiljer sig från fallet med statliga stöd som beviljats i strid med gällande rätt. De senare kan enligt rättspraxis inte ”läkas” i efterhand. I förevarande mål rör frågan gränserna för en medlemsstats unionsrättsliga skyldigheter snarare än följderna av en överträdelse av dessa. Se dom av den 21 oktober 2003 i de förenade målen C-261/01 och C-262/01, van Calster m.fl. (REG 2003, s. I-12249).
Dom av den 13 mars 2007 i mål C-524/04,Test Claimants in the Thin Cap Group Litigation (REG 2007, s. I-2107), punkterna 98–100.
Det ska påpekas att section 402(3A) och (3B) ICTA, vilka infördes år 2000, föregicks av en bestämmelse enligt vilken ”bolag” endast avsåg bolag i Förenade kungariket. Se section 258(7) ICTA 1970 (återgiven i domen i det ovannämnda målet ICI, punkt 6).
Såsom generaladvokaten har angett i punkterna 182–184 i sitt förslag till avgörande begränsar de villkor som ställs i direktiv 96/61 äganderätten när det gäller områden som berörs av en anläggning som omfattas av direktivets tillämpningsområde.
Äganderätten ska emellertid inte betraktas som en absolut rättighet, utan måste bedömas utifrån sin funktion i samhället. Följaktligen kan begränsningar införas i utövandet av äganderätten, förutsatt att begränsningarna verkligen svarar mot mål av allmänintresse och inte innebär ett, i förhållande till det eftersträvade målet, orimligt och icke godtagbart ingrepp som påverkar kärnan i denna rättighet (dom av den 3 september 2008 i de förenade målen C-402/05 P och C-415/05 P, Kadi och Al Barakaat International Foundation mot rådet och kommissionen, REG 2008, s. I-6351, punkt 355 och av den 9 mars 2010 i de förenade målen C-379/08 och C-380/08, ERG m.fl., REU 2010, s. I-2007, punkt 80).
Vad avser de mål av allmänintresse som nämnts ovan framgår det av fast rättspraxis att miljöskydd ingår bland dessa mål och således kan motivera en begränsning av utövandet av äganderätten (se dom av den 7 februari 1985 i mål 240/83, ADBHU, REG 1985, s. 531, punkt 13, av den 20 september 1988 i mål 302/86, kommissionen mot Danmark, REG 1988, s. 4607, punkt 8, svensk specialutgåva, volym 9, s. 579, av den 2 april 1998 i mål C-213/96, Outokumpu, REG 1998, s. I-1777, punkt 32, och domen i de ovannämnda förenade målen ERG m.fl., punkt 81).
När det gäller frågan huruvida det aktuella ingreppet i äganderätten, för det fall det visar sig föreligga ett sådant, är proportionerligt räcker det att konstatera att direktiv 96/61 upprätthåller en balans mellan de krav som är knutna till äganderätten och miljöskyddskraven.
Mot denna bakgrund ska den femte frågan besvaras enligt följande: Ett avgörande från en nationell domstol, som fattats inom ramen för ett nationellt förfarande genom vilket medlemsstaten uppfyller sina åtaganden enligt artikel 15a i direktiv 96/91 och artikel 9.2 och 9.4 i Århuskonventionen och som upphäver ett tillstånd som beviljats i strid med bestämmelserna i nämnda direktiv, kan inte som sådant utgöra ett oberättigat ingrepp i exploatörens äganderätt enligt artikel 17 i Europeiska unionens stadga om de grundläggande rättigheterna.
Rättegångskostnader
Eftersom förfarandet i förhållande till parterna i målet vid den nationella domstolen utgör ett led i beredningen av samma mål, ankommer det på den nationella domstolen att besluta om rättegångskostnaderna. De kostnader för att avge yttranden till domstolen som andra än nämnda parter har haft är inte ersättningsgilla.
Mot denna bakgrund beslutar domstolen (stora avdelningen) följande:
Artikel 267 FEUF ska tolkas så, att en nationell domstol, såsom den hänskjutande domstolen, är skyldig att på eget initiativ begära förhandsavgörande från Europeiska unionens domstol även om det mål den har att avgöra har återförvisats till den efter det att dess första avgörande i saken upphävts av författningsdomstolen i den aktuella medlemsstaten och den, enligt en nationell bestämmelse, är skyldig att lägga författningsdomstolens rättsliga bedömning till grund för sitt avgörande av tvisten.
Rådets direktiv 96/61/EG av den 24 september 1996 om samordnade åtgärder för att förebygga och begränsa föroreningar, i dess lydelse enligt Europaparlamentets och rådets förordning (EG) nr 166/2006 av den 18 januari 2006, ska tolkas så, att det
kräver att den berörda allmänheten ges tillgång till ett stadsplaneringsbeslut, såsom det som är i fråga i det nationella målet, redan från det att tillståndsförfarandet avseende den aktuella anläggningen inleds,
inte tillåter att de behöriga nationella myndigheterna nekar den berörda allmänheten tillgång till ett sådant beslut med hänvisning till skyddet för sekretess som omfattar kommersiell eller industriell information, där sådan sekretess föreskrivs i nationell lagstiftning eller unionslagstiftning i syfte att skydda legitima ekonomiska intressen, och
inte utgör hinder för att en oberättigad vägran att ge den berörda allmänheten tillgång till ett sådant stadsplaneringsbeslut som det nationella målet avser under det administrativa förfarandet i första instans kan rättas till under det administrativa förfarandet i andra instans, under förutsättning att alla alternativ fortfarande är möjliga och att en rättelse i detta skede i förfarandet innebär att allmänheten fortfarande kan delta på ett meningsfullt sätt i beslutsförfarandet. Det ankommer på den nationella domstolen att pröva huruvida så är fallet.
Artikel 15a i direktiv 96/61, i dess lydelse enligt förordning nr 166/2006, ska tolkas så, att medlemmarna av den berörda allmänheten, inom ramen för en sådan rättslig prövning som föreskrivs i denna bestämmelse, ska ha rätt att yrka att den domstol eller annat oberoende och opartiskt behörigt organ som inrättats genom lag ska förordna om interimistiska åtgärder i form av inhibition av ett tillstånd enligt artikel 4 i direktivet intill dess att ett slutligt avgörande meddelas.
Ett avgörande från en nationell domstol, som fattats inom ramen för ett nationellt förfarande genom vilket medlemsstaten uppfyller sina åtaganden enligt artikel 15a i direktiv 96/91, i dess lydelse enligt förordning nr 166/2006, och artikel 9.2 och 9.4 i konventionen om tillgång till information, allmänhetens deltagande i beslutsprocesser och tillgång till rättslig prövning i miljöfrågor, som undertecknades i Århus den 25 juni 1998 och som godkändes på Europeiska gemenskapens vägnar genom rådets beslut 2005/370/EG av den 17 februari 2005, och som upphäver ett tillstånd som beviljats i strid med bestämmelserna i nämnda direktiv, kan inte som sådant utgöra ett oberättigat ingrepp i exploatörens äganderätt enligt artikel 17 i Europeiska unionens stadga om de grundläggande rättigheterna.
Begäran om förhandsavgörande — Område med frihet, säkerhet och rättvisa — Direktiv 2004/83/EG — Miniminormer för beviljande av flyktingstatus eller status som alternativt skyddsbehövande — Artikel 4 — Bedömning av fakta och omständigheter — Bedömningsmetoder — Godtagande av viss bevisning — Omfattningen av de behöriga nationella myndigheternas befogenheter — Fruktan för förföljelse på grund av sexuell läggning — Skillnader mellan å ena sidan gränserna för bedömningen av uppgifter och skriftliga eller andra bevis avseende en asylsökandes påstådda sexuella läggning och å andra sidan motsvarande gränser avseende andra skäl för förföljelse — Direktiv 2005/85/EG — Miniminormer för medlemsstaternas förfaranden för beviljande eller återkallande av flyktingstatus — Artikel 13 — Krav på den personliga intervjun — Europeiska unionens stadga om de grundläggande rättigheterna — Artikel 1 — Människans värdighet — Artikel 7 — Respekt för privatlivet och familjelivet”
I de förenade målen C‑148/13–C‑150/13,
angående tre beslut att begära förhandsavgörande enligt artikel 267 FEUF, från Raad van State (Nederländerna), av den 20 mars 2013, som inkom till domstolen den 25 mars 2013, i målen
A (C‑148/13),
B (C‑149/13),
C (C‑150/13)
mot
Staatssecretaris van Veiligheid en Justitie,
ytterligare deltagare i rättegången:
United Nations High Commissioner for Refugees (UNHCR),
meddelar
DOMSTOLEN (stora avdelningen)
sammansatt av ordföranden V. Skouris, vice-ordföranden K. Lenaerts, avdelningsordförandena A. Tizzano, L. Bay Larsen (referent), T. von Danwitz, A. Ó Caoimh och J.-C. Bonichot, samt domarna A. Borg Barthet, J. Malenovský, E. Levits, E. Jarašiūnas, C.G. Fernlund och J.L. da Cruz Vilaça,
generaladvokat: E. Sharpston,
justitiesekreterare: förste handläggaren M. Ferreira,
efter det skriftliga förfarandet och förhandlingen den 25 februari 2014,
med beaktande av de yttranden som avgetts av:
A, genom N.C. Blomjous, advocaat,
B, genom C. Chen, advocaat,
United Nations High Commissioner for Refugees (UNHCR), genom P. Moreau, i egenskap av ombud, biträdd av M.-E. Demetriou, QC,
Nederländernas regering, genom C. Schillemans, M. Bulterman och B. Koopman, samtliga i egenskap av ombud,
Belgiens regering, genom M. Jacobs och C. Pochet, båda i egenskap av ombud,
Tjeckiens regering, genom M. Smolek och J. Vláčil, båda i egenskap av ombud,
Tysklands regering, genom T. Henze och A. Wiedmann, båda i egenskap av ombud,
Greklands regering, genom M. Michelogiannaki, i egenskap av ombud,
Frankrikes regering, genom D. Colas och S. Menez, båda i egenskap av ombud,
Europeiska kommissionen, genom M. Condou-Durande och R. Troosters, båda i egenskap av ombud,
och efter att den 17 juli 2014 ha hört generaladvokatens förslag till avgörande,
följande
Dom
Respektive begäran om förhandsavgörande avser tolkningen av artikel 4 i rådets direktiv 2004/83/EG av den 29 april 2004 om miniminormer för när tredjelandsmedborgare eller statslösa personer skall betraktas som flyktingar eller som personer som av andra skäl behöver internationellt skydd samt om dessa personers rättsliga ställning och om innehållet i det beviljade skyddet (EUT L 304, s. 12, med rättelse i EUT L 204, 2005, s. 24, och i EUT L 278, 2011, s. 13), samt av artiklarna 3 och 7 i Europeiska unionens stadga om de grundläggande rättigheterna (nedan kallad stadgan).
Respektive begäran har framställts i mål mellan å ena sidan tredjelandsmedborgarna A, B respektive C, och å andra sidan Staatssecretaris van Veiligheid en Justitie (statssekreteraren för säkerhetsfrågor och justitiefrågor) (nedan kallad Staatssecretaris). Målen rör nämnda tredjelandsmedborgares ansökningar om tillfälligt uppehållstillstånd (asyl) i Nederländerna.
Tillämpliga bestämmelser
Internationell rätt
Konventionen angående flyktingars rättsliga ställning undertecknades i Genève den 28 juli 1951 (Förenta nationernas fördragssamling, volym 189, s. 150, nr 2545 (1954)) och trädde i kraft den 22 april 1954. Den har kompletterats genom protokollet angående flyktingars rättsliga ställning, som antogs i New York den 31 januari 1967 och trädde i kraft den 4 oktober 1967 (nedan kallad Genèvekonventionen). I artikel 1 A punkt 2 första stycket i Genèvekonventionen föreskrivs att med uttrycket ”flykting”avses den som ”i anledning av välgrundad fruktan för förföljelse på grund av sin ras, religion, nationalitet, tillhörighet till viss samhällsgrupp eller politiska åskådning befinner sig utanför det land, vari han är medborgare, samt är ur stånd att eller på grund av sådan fruktan, som nyss sagts, icke önskar att begagna sig av sagda lands skydd eller den som, utan att vara medborgare i något land, till följd av händelser som förut sagts befinner sig utanför det land, vari han tidigare haft sin vanliga vistelseort, samt är ur stånd att eller på grund av sådan fruktan, som nyss sagts, icke önskar att återvända dit”.
Unionsrätt
Direktiv 2004/83
Enligt skäl 3 i direktiv 2004/83 utgör Genèvekonventionen grundstenen i det folkrättsliga systemet för skydd av flyktingar.
I skäl 10 i direktivet anges följande:
Detta direktiv står i överensstämmelse med de grundläggande rättigheter och principer som erkänns särskilt i [stadgan]. Direktivet syftar särskilt till att säkerställa full respekt för den mänskliga värdigheten och de asylsökandes och deras medföljande familjemedlemmars rätt till asyl.”
I skäl 16 i direktivet anges att det bör fastställas miniminormer för definitionen och innebörden av flyktingstatus för att vägleda medlemsstaternas behöriga myndigheter vid tillämpningen av Genèvekonventionen.
Enligt skäl 17 i direktiv 2004/83 är det nödvändigt att införa gemensamma kriterier för när asylsökande ska erkännas som flyktingar i den mening som avses i artikel 1 i Genèvekonventionen.
Det anges i artikel 2 i direktivet att följande beteckningar används i det direktivet med de betydelser som här anges:
...
’flykting’, en tredjelandsmedborgare som med anledning av välgrundad fruktan för förföljelse på grund av ras, religion, nationalitet, politisk åskådning eller tillhörighet till viss samhällsgrupp befinner sig utanför det land där han eller hon är medborgare och som inte kan eller på grund av sin fruktan inte vill begagna sig av det landets skydd …
...”
I artikel 4 i direktiv 2004/83, som återfinns i direktivets kapitel II med rubriken ”Bedömning av ansökningar om internationellt skydd”, uppställs villkoren för bedömningen av fakta och omständigheter. Där anges följande:
1.   Medlemsstaterna får betrakta det som den sökandes skyldighet att så snart som möjligt lägga fram alla faktorer som behövs för att styrka ansökan om internationellt skydd. Det är medlemsstaternas skyldighet att i samarbete med den sökande bedöma de relevanta faktorerna i ansökan.
De faktorer som det hänvisas till i punkt 1 utgörs av den sökandes utsagor och alla handlingar som den sökande förfogar över angående den sökandes ålder, bakgrund, inklusive relevanta släktingars bakgrund, identitet, nationalitet(er), tidigare bosättningsland(länder) och -ort(er), tidigare asylansökningar, resvägar, identitets- och resehandlingar samt orsakerna till ansökan om internationellt skydd.
Bedömningen av en ansökan om internationellt skydd skall vara individuell, och följande skall beaktas:
Alla relevanta uppgifter om ursprungslandet vid den tidpunkt då beslut fattas om ansökan, inbegripet lagar och andra författningar i ursprungslandet samt det sätt på vilket dessa tillämpas.
De relevanta utsagor och handlingar som den sökande har lämnat, inklusive information om huruvida sökanden har varit eller kan bli utsatt för förföljelse eller allvarlig skada.
Sökandens personliga ställning och förhållanden, inklusive faktorer som bakgrund, kön och ålder, så att det kan bedömas huruvida de handlingar den sökande har blivit eller skulle kunna bli utsatt för, på grundval av sökandens personliga omständigheter, skulle innebära förföljelse eller allvarlig skada.
Om den sökande efter att ha lämnat ursprungslandet ägnat sig åt en verksamhet, vars enda syfte eller vars huvudsyfte var att skapa de nödvändiga förutsättningarna för att ansöka om internationellt skydd, skall man bedöma om denna verksamhet kommer att utsätta den sökande för förföljelse eller allvarlig skada om han eller hon återvänder till landet.
Om man rimligen kan förvänta sig att den sökande begagnar sig av skyddet i ett annat land där han eller hon kan hävda sitt medborgarskap.
...
När medlemsstaterna tillämpar principen enligt vilken det är den sökandes skyldighet att styrka sin ansökan om internationellt skydd, och den sökandes uppgifter inte kan styrkas av skriftliga eller andra bevis, skall sådana uppgifter inte behöva bekräftas om följande villkor är uppfyllda:
Sökanden har gjort en genuin ansträngning för att styrka sin ansökan.
Alla relevanta faktorer som den sökande förfogar över har lagts fram och en tillfredsställande förklaring har lämnats till varför andra relevanta faktorer saknas.
Sökandens uppgifter befinns vara sammanhängande och rimliga och strider inte mot tillgänglig specifik och allmän information som rör den sökandes ärende.
Sökanden har ansökt om internationellt skydd så tidigt som möjligt, såvida inte sökanden kan framföra goda skäl till varför han eller hon inte gjort det.
Sökandens allmänna trovärdighet är fastställd.”
Artikel 10 i direktiv 2004/83, med rubriken ”Skäl till förföljelsen”, innehåller följande bestämmelser:
1.   Medlemsstaterna skall ta hänsyn till följande faktorer vid bedömningen av skälen till förföljelsen:
...
En grupp skall anses utgöra en särskild samhällsgrupp, särskilt när
gruppens medlemmar har en gemensam väsentlig egenskap eller en gemensam bakgrund som inte kan ändras, eller består av personer som har en gemensam egenskap eller övertygelse som är så grundläggande för identiteten eller samvetet att de inte får tvingas avsvära sig den,
gruppen har en särskild identitet i det berörda landet eftersom den uppfattas som annorlunda av omgivningen.
Beroende på omständigheterna i ursprungslandet kan en särskild samhällsgrupp omfatta en grupp grundad på en gemensam egenskap, till exempel sexuell läggning. Sexuell läggning får inte tolkas så att det innefattar handlingar som anses brottsliga enligt medlemsstaternas nationella lagstiftning. ...
...”
Direktiv 2005/85/EG
I skäl 8 i rådets direktiv 2005/85/EG av den 1 december 2005 om miniminormer för medlemsstaternas förfaranden för beviljande eller återkallande av flyktingstatus (EUT L 326, s. 13, och rättelse i EUT L 236, 2006, s. 36) anges att detta direktiv står i överensstämmelse med de grundläggande rättigheter och principer som erkänns särskilt i Europeiska unionens stadga om de grundläggande rättigheterna.
I artikel 13 i direktiv 2005/85 preciseras kraven på den personliga intervjun och i punkt 3 föreskrivs följande:
Medlemsstaterna skall vidta lämpliga åtgärder för att se till att personliga intervjuer genomförs under sådana förhållanden att sökandena kan lägga fram skälen för sina ansökningar på ett heltäckande sätt. Medlemsstaterna skall därför:
se till att intervjuaren är tillräckligt kompetent för att om möjligt kunna beakta de personliga och allmänna omständigheter som ligger bakom ansökan, inklusive sökandens kulturella ursprung eller utsatta ställning …
...”
Nederländsk rätt
Den relevanta nederländska lagstiftningen återfinns i artikel 31 i 2000 års utlänningslag (Vreemdelingenwet 2000), artikel 3.111 i 2000 års utlänningsförordning (Vreemdelingenbesluit 2000) och artikel 3.35 i 2000 års utlänningsföreskrifter (Voorschrift Vreemdelingen 2000).
Riktlinjer om hur dessa bestämmelser ska tolkas finns i 2000 års utlänningscirkulär (Vreemdelingencirculaire 2000), punkterna C2/2.1, C2/2.1.1 och C14/2.1–C14/2.4.
Det framgår av artikel 31.1 i 2000 års utlänningslag, jämförd med artikel 3.111 punkt 1 i 2000 års utlänningsförordning, att det ankommer på den asylsökande att göra de uppgifter som har åberopats till stöd för ansökan om tillfälligt uppehållstillstånd (asyl) sannolika och att vederbörande är skyldig att på eget initiativ tillhandahålla samtliga relevanta uppgifter som myndigheten behöver för att kunna fatta beslut i ärendet. Staatssecretaris gör en bedömning av huruvida det finns stöd i lag för att bevilja ett sådant uppehållstillstånd.
Det framgår av artikel 3.111 punkt 1 i 2000 års utlänningsförordning att när en asylsökande ansöker om ett sådant uppehållstillstånd som avses i artikel 28 i 2000 års utlänningslag, ska han eller hon tillhandahålla samtliga uppgifter, inklusive relevanta handlingar, som Staatssecretaris kan lägga till grund för den bedömning av huruvida det föreligger rättsligt stöd för ett bifall av ansökan som görs i samarbete med asylsökanden.
Enligt punkt C14/2.1 i 2000 års utlänningscirkulär ska bedömningen av trovärdigheten i de uppgifter som en asylsökande har lämnat omfatta de fakta och omständigheter som han eller hon har gjort gällande. De faktiska omständigheterna är uppgifter som rör den asylsökandes person, bland annat personens sexuella läggning.
I punkt C14/2.2 i cirkuläret anges att en asylsökande är skyldig att säga sanningen och att fullt ut samarbeta för att bidra till att samtliga omständigheter kan klarläggas på ett så fullständigt sätt som möjligt. Vederbörande är skyldig att så snart som möjligt informera myndigheten för immigrations- och medborgarskapsfrågor om alla händelser och faktiska omständigheter som är av betydelse för handläggningen av ärendet.
Det anges i punkt C14/2.3 i cirkuläret att om en del av en asylsökandes berättelse brister i trovärdighet är det inte uteslutet att detta även sänker berättelsens trovärdighet i övriga delar.
Det framgår av punkt C14/2.4 i cirkuläret att det i princip räcker med att en asylsökande har gjort sin berättelse sannolik. För detta förväntas vederbörande inkomma med handlingar till stöd för sin ansökan. Trovärdighetsbedömningen av de uppgifter som den asylsökande har lämnat till stöd för sin ansökan handlar emellertid inte om huruvida, och i så fall i vilken utsträckning, dessa uppgifter kan styrkas. I många fall har nämligen asylsökande visat att de saknar möjlighet att styrka sina uppgifter och att det inte rimligen kan krävas att de inger övertygande bevisning till stöd för sina berättelser.
Staatssecretaris har möjlighet att betrakta uppgifterna som trovärdiga med stöd av artikel 3.35 punkt 3 i 2000 års utlänningsföreskrifter och således inte kräva någon bekräftelse av dessa om den asylsökandes allmänna trovärdighet har kunnat fastställas.
Målen vid den nationella domstolen och tolkningsfrågan
Tredjelandsmedborgarna A, B och C ingav varsin ansökan om tillfälligt uppehållstillstånd (asyl) i Nederländerna. Till stöd för sina ansökningar gjorde de gällande att de fruktade förföljelse i sina respektive ursprungsländer, framför allt på grund av deras homosexuella läggning.
Den första asylansökan, som hade ingetts av A, avslogs av Staatssecretaris med hänvisning till bristande trovärdighet.
A bestred inte detta första avslagsbeslut. I stället inkom han med en andra asylansökan, varvid han uppgav sig vara beredd att genomgå ett ”test” som skulle styrka hans homosexuella läggning eller att utföra en sexuell handling för att bevisa att hans sexuella läggning var den han påstod.
Staatssecretaris beslutade den 12 juli 2011 att avslå A:s andra ansökan med motiveringen att vederbörandes påstående om sexuell läggning fortfarande inte var trovärdigt. Staatssecretaris fann att man inte kunde godta påståendet om den asylsökandes sexuella läggning utan att göra någon bedömning av sökandens trovärdighet.
Den 1 augusti 2012 avslog Staatssecretaris B:s ansökan med motiveringen att den redogörelse som lämnats beträffande B:s homosexuella läggning var vag, knapphändig och inte trovärdig. Dessutom fann Staatssecretaris att eftersom B kom från ett land där homosexualitet inte är accepterat borde vederbörande ha kunnat redogöra mer i detalj för sina känslor och för den inre process som han genomgått vad gäller sin sexuella läggning.
C ingav en första asylansökan. Till stöd för ansökan åberopade han andra grunder än förföljelse på grund av homosexualitet. Ansökan avslogs av Staatssecretaris.
C bestred inte detta första avslagsbeslut. Istället inkom han med en andra asylansökan, denna gång med åberopande av att han kände fruktan för förföljelse i ursprungslandet på grund av sin homosexuella läggning. I samband med denna andra ansökan hävdade C att han inte hade insett att han var homosexuell förrän efter det att han hade lämnat sitt ursprungsland. Till stöd för sin ansökan gav C till de myndigheter som ansvarade för handläggningen av hans ärende in en videoupptagning som visar intima handlingar som utförs tillsammans med en person av samma kön.
Den 8 oktober 2012 avslog Staatssecretaris C:s asylansökan med motiveringen att hans redogörelser för sin homosexuella läggning inte var trovärdiga. Staatssecretaris fann att C borde ha nämnt sin homosexuella läggning i samband med sin första asylansökan, att C inte hade lämnat någon tydlig förklaring till hur han hade blivit medveten om sin homosexuella läggning och att han inte hade kunnat svara på frågor om nederländska organisationer som försvarar homosexuellas rättigheter.
A, B och C överklagade besluten att avslå deras ansökningar om tillfälligt uppehållstillstånd (asyl) till Rechtbank ’s-Gravenhage (nedan kallad Rechtbank).
Rechtbank ogillade A:s och C:s överklaganden genom domar som meddelades den 9 september 2011 och den 30 oktober 2012. Rechtbank fann för det första att A och C i sina överklaganden borde ha bestritt de första avslagsbesluten från Staatssecretaris, och för det andra att de inte under det andra asylförfarandet hade lyckats göra sina redogörelser för den påstådda homosexuella läggningen trovärdiga.
Genom dom av den 23 augusti 2012 ogillade Rechtbank likaså B:s överklagande av Staatssecretaris avslagsbeslut. Rechtbank bedömde att Staatssecretaris hade haft rimligt fog för slutsatsen att B:s redogörelse för sin homosexuella läggning inte var trovärdig.
A, B och C överklagade domarna till Raad van State.
I målen om överklagande har A, B och C framför allt gjort gällande att det är omöjligt att objektivt fastställa en asylsökandes sexuella läggning. När de myndigheter som prövar en asylansökan fattar sitt beslut måste de därför godta en asylsökandes påstående som sådant vad gäller hans eller hennes sexuella läggning.
A, B och C har emellertid gjort gällande att dessa myndigheter, vid bedömningen av trovärdigheten i de uppgifter som den asylsökande har lämnat, ställer frågor om den påstådda läggningen, vilka är av sådan art att de inkräktar på bland annat den asylsökandes värdighet och hans eller hennes rätt till respekt för privatlivet. Dessutom tas ingen hänsyn till det obehag som den asylsökande kan uppleva under förhören eller till de kulturella barriärer som kan hindra honom eller henne från att tala öppet om sin läggning. Därtill anser A, B och C att det faktum att Staatssecretaris finner att en asylberättelse framstår som inte trovärdig inte får leda till att samma slutsats dras vad gäller trovärdighetsbedömningen av den sexuella läggningen i sig.
Staatssecretaris har påpekat att det inte framgår av vare sig direktiv 2004/83 eller av stadgan att beslut ska fattas på grundval enbart av de asylsökandes påstående om sexuell läggning. Det som ska kontrolleras är emellertid inte huruvida de asylsökande verkligen har den sexuella läggning som de påstår sig ha, utan huruvida de har gjort det sannolikt att de tillhör en samhällsgrupp i den mening som avses i artikel 10.1 d i direktiv 2004/83 eller att de som utövar förföljelse betraktar dem som sådana i den mening som avses i artikel 10.2 i direktivet.
Dessutom har Staatssecretaris konstaterat att det är mycket sällsynt att en asylsökande kan bevisa sin homosexuella läggning annat än genom sin egen berättelse, vilket betyder att när denna berättelse anses vara sammanhängande och sannolik och det har kunnat fastställas att den asylsökande är allmänt trovärdig ska vederbörande tillerkännas förmånen av uppkommet tvivelsmål.
Enligt Staatssecretaris skiljer sig den trovärdighetsbedömning som ska göras beträffande asylsökandes sexuella läggning inte från den som ska göras när det är andra skäl för förföljelse som åberopas. Denna myndighet tar dock hänsyn till att uppgifter om sexuell läggning är förenade med särskilda problem. Bland annat rekommenderas de medarbetare som sköter intervjuerna med de asylsökande att inte ställa direkta frågor om på vilket sätt de asylsökande lever ut sin läggning. Dessutom har Staatssecretaris uppgett att bilder av intima handlingar som har lämnats in som bevisning av de asylsökande inte tillmäts någon betydelse, eftersom dessa bilder endast styrker utförandet i sig av sexuella handlingar och inte den påstådda sexuella läggningen i sig.
Raad van State har förtydligat att varken artikel 4 i direktiv 2004/83 eller de åberopade bestämmelserna i stadgan innehåller någon skyldighet för Staatssecretaris att godta de asylsökandes påståenden som sådana för att betrakta deras sexuella läggning som styrkt. Dessutom konstaterar Raad van State att prövningen av asylsökandes sexuella läggning inte skiljer sig från prövningen av andra skäl till förföljelse.
Raad van State undrar dock om det genom bestämmelserna i artikel 4 i direktiv 2004/83 och bestämmelserna i artiklarna 3 och 7 i stadgan uppställs några eventuella gränser för hur bedömningen av de asylsökandes sexuella läggning får göras.
Att ställa frågor till den asylsökande kan enligt Raad van State i viss mån inkräkta på de rättigheter som garanteras genom de ovannämnda bestämmelserna i stadgan.
Raad van State anser att det oavsett vilken metod som den berörda medlemsstaten har valt för att bedöma sanningshalten i ett påstående om sexuell läggning inte kan uteslutas att det finns en risk för att inkräkta på de asylsökandes grundläggande rättigheter enligt artiklarna 3 och 7 i stadgan.
Mot denna bakgrund beslutade Raad van State att vilandeförklara målet och att till domstolen hänskjuta följande fråga, vilken har formulerats på samma sätt i vart och ett av målen C‑148/13–C‑150/13:
Vilka gränser för sättet att genomföra en trovärdighetsbedömning av ett påstående om viss sexuell läggning uppställs genom artikel 4 i [direktiv 2004/83] och genom [stadgan], framför allt artiklarna 3 och 7, och skiljer sig dessa gränser från dem som gäller för trovärdighetsbedömningen av andra skäl till förföljelse, och i så fall i vilket avseende?”
Domstolen beslutade den 19 april 2013 att förena målen C‑148/13–C‑150/13 vad gäller det skriftliga och det muntliga förfarandet samt domen.
Prövning av tolkningsfrågan
Inledande synpunkter
Det framgår av skälen 3, 16 och 17 i direktiv 2004/83 att Genèvekonventionen utgör grundstenen i det folkrättsliga systemet för skydd av flyktingar och att bestämmelserna i direktivet om villkoren för beviljande av flyktingstatus och om innebörden av flyktingstatus har antagits för att hjälpa medlemsstaternas behöriga myndigheter att tillämpa Genèvekonventionen på grundval av gemensamma begrepp och kriterier (dom N., C‑604/12, EU:C:2014:302, punkt 27).
Bestämmelserna i direktiv 2004/83 ska således tolkas mot bakgrund av direktivets systematik och syfte, med beaktande av Genèvekonventionen och de andra relevanta fördrag som avses i artikel 78.1 FEUF. Såsom framgår av skäl 10 i direktivet ska tolkningen även stå i överensstämmelse med de rättigheter som erkänns i stadgan (dom X m.fl., C‑199/12–C‑201/12, EU:C:2013:720, punkt 40).
Vidare ska det erinras om att direktiv 2004/83 inte innehåller några förfaranderegler för prövningen av en ansökan om internationellt skydd och således inte heller några rättssäkerhetsgarantier för den asylsökande. Det är i direktiv 2005/85 som det fastställs miniminormer för förfarandena vid prövningen av ansökningar, och det är även i det direktivet som man återfinner bestämmelserna om de asylsökandes rättigheter, vilka ska beaktas vid prövningen av de nu aktuella nationella målen.
Frågan
Den hänskjutande domstolen har ställt sin fråga för att få klarhet i huruvida artikel 4 i direktiv 2004/83, jämförd med bestämmelserna i stadgan, ska tolkas så, att den uppställer vissa gränser för den bedömning av fakta och omständigheter som de behöriga nationella myndigheterna får göra – och som kan bli föremål för prövning i domstol – för att fastställa den sexuella läggningen hos en asylsökande, som till stöd för sin asylansökan har åberopat fruktan för förföljelse på grund av denna läggning.
I det avseendet har A, B och C hävdat att de behöriga myndigheter som har i uppgift att pröva en asylansökan till stöd för vilken den asylsökande har åberopat fruktan för förföljelse på grund av sexuell läggning måste godta den påstådda läggningen som en styrkt omständighet redan på grundval av den asylsökandes uppgifter. Domstolen finner dock, med hänsyn till asylförfarandets särskilda sammanhang, att dessa uppgifter inte kan utgöra något annat än utgångspunkten i processen för att bedöma fakta och omständigheter enligt artikel 4 i direktiv 2004/83.
Det framgår nämligen av själva lydelsen i artikel 4.1 i direktivet att medlemsstaterna får betrakta det som den sökandes skyldighet att så snart som möjligt lägga fram alla faktorer som behövs för att styrka ansökan om internationellt skydd och att det är deras skyldighet att i samarbete med den sökande bedöma de relevanta faktorerna i ansökan.
Dessutom följer det av artikel 4.5 i direktiv 2004/83 att när villkoren i punkterna a–e inte är uppfyllda, kan asylsökandes uppgifter om deras påstådda sexuella läggning behöva bekräftas.
Således konstaterar domstolen att även om det ankommer på den asylsökande att informera om sin läggning, vilken utgör en personlig angelägenhet, kan asylansökningar till stöd för vilka sökanden har åberopat en fruktan för förföljelse på grund av denna läggning, precis som de ansökningar som grundas på andra skäl för förföljelse, bli föremål för en bedömningsprocess enligt artikel 4 i direktivet.
Dock måste de metoder som de behöriga myndigheterna använder för att bedöma de uppgifter och skriftliga eller andra bevis som har åberopats till stöd för sådana ansökningar vara förenliga med bestämmelserna i direktiven 2004/83 och 2005/85 och även – såsom framgår av skäl 10 respektive skäl 8 i dessa direktiv – med de grundläggande rättigheter som garanteras genom stadgan, såsom rätten till människans värdighet (artikel 1 i stadgan) och rätten till respekt för privatlivet och familjelivet (artikel 7 i stadgan).
Visserligen är bestämmelserna i artikel 4 i direktiv 2004/83 tillämpliga på samtliga ansökningar om internationellt skydd, oavsett vilka skäl för förföljelse som har åberopats till stöd för dessa. Det hindrar emellertid inte att det ankommer på de behöriga myndigheterna att anpassa de metoder som används vid bedömningen av uppgifter och skriftliga eller andra bevis utifrån vad som kännetecknar olika typer av asylansökningar, och att iaktta de rättigheter som garanteras genom stadgan.
Såsom domstolen konstaterade i punkt 64 i domen M (C‑277/11, EU:C:2012:744) kan ska bedömningen av fakta och omständigheter enligt artikel 4 i direktiv 2004/83 göras i två led. Först ska det fastställas vilka faktiska omständigheter som kan utgöra bevis till stöd för ansökan. Därefter ska det göras en rättslig prövning av dessa omständigheter. Under den rättsliga prövningen ska det mot bakgrund av omständigheterna i det enskilda fallet avgöras huruvida de materiella förutsättningar för att beviljas internationellt skydd som föreskrivs i artiklarna 9 och 10 eller 15 i direktiv 2004/83 är uppfyllda.
När det gäller det första skedet, som Raad van States frågor i samtliga av de nationella målen just handlar om, finner domstolen att även om medlemsstaterna normalt sett får betrakta det som en skyldighet för den sökande – vilken för övrigt är den som är bäst lämpad för att lämna uppgifter till stöd för den egna sexuella läggningen – att lägga fram alla faktorer som behövs för att styrka ansökan, är den berörda medlemsstaten dock skyldig att samarbeta med den sökande vid fastställandet av de för ansökan relevanta faktorerna i enlighet med artikel 4.1 i direktivet (se, för ett liknande resonemang, dom M., EU:C:2012:744, punkt 65).
Enligt artikel 4.3 c i direktiv 2004/83 ska denna bedömning vara individuell och göras med beaktande av sökandens personliga ställning och förhållanden, inklusive faktorer som bakgrund, kön och ålder, så att det kan bedömas huruvida de handlingar den sökande har blivit eller skulle kunna bli utsatt för, på grundval av dessa personliga förhållanden, skulle innebära förföljelse eller allvarlig skada.
Härtill kommer, såsom det erinras om ovan i punkt 51, att det i artikel 4 i nämnda direktiv anges att när en asylsökandes uppgifter inte kan styrkas av skriftliga eller andra bevis, ska sådana uppgifter, vid de behöriga myndigheternas bedömning, inte behöva bekräftas om de kumulativa villkoren i artikel 4.5 a–e i direktivet är uppfyllda.
Domstolen övergår därefter till att behandla metoderna för att bedöma de uppgifter och skriftliga eller andra bevis som är i fråga i vart och ett av de nationella målen. För att Raad van State ska få ett användbart svar kommer prövningen att begränsas till två frågeställningar. För det första ska det prövas huruvida det är förenligt med bestämmelserna i direktiven 2004/83 och 2005/85 samt bestämmelserna i stadgan dels att de behöriga myndigheterna genomför kontroller med hjälp av förhör baserade på bland annat stereotyper av homosexuella eller detaljerade förhör om den asylsökandes sexuella vanor, dels att dessa myndigheter kan godta att den asylsökande genomgår ”test” för fastställande av personens homosexuella läggning och/eller, på frivillig basis, ge in videoupptagningar som visar när vederbörande utför intima handlingar. För det andra ska det prövas huruvida det är förenligt med ovannämnda bestämmelser att de behöriga myndigheterna redan av det skälet att den asylsökande inte åberopade sin påstådda sexuella läggning första gången han eller hon gavs tillfälle att lägga fram skälen till förföljelse kan dra slutsatsen att den asylsökande brister i trovärdighet.
När det gäller bedömningar som grundas på förhör om den asylsökandes kunskaper om sådana organisationer som tillvaratar homosexuellas intressen och om detaljer beträffande dessa, har klaganden i det nationella målet i mål C‑150/13 hävdat att sådana förhör innebär att myndigheterna grundar sina bedömningar på stereotypa uppfattningar om homosexuellas beteenden och inte på den konkreta situation som den enskilda asylsökanden befinner sig i.
I det avseendet föreskrivs, som redan angetts, i artikel 4.3 c i direktiv 2004/83 att de behöriga myndigheterna ska göra sin bedömning med beaktande av sökandens personliga ställning och förhållanden och i artikel 13.3 a i direktiv 2005/85 att dessa myndigheter vid en intervju ska beakta de personliga och allmänna omständigheter som ligger bakom ansökan.
Visserligen kan förhör som grundas på stereotypa uppfattningar vara användbara för de behöriga myndigheterna när de gör sin bedömning. En asylprövning som uteslutande baseras på stereotypa uppfattningar om homosexuella uppfyller dock inte kraven i de bestämmelser som avses i föregående punkt, eftersom nämnda myndigheter då inte ges möjlighet att beakta den asylsökandes individuella och personliga förhållanden.
En asylsökandes oförmåga att svara på sådana frågor räcker således inte i sig som skäl för att slå fast att vederbörande brister i trovärdighet, eftersom ett sådant tillvägagångssätt skulle strida mot kraven i artikel 4.3 c i direktiv 2004/83 och artikel 13.3 a i direktiv 2005/85.
Vidare konstaterar domstolen att även om de nationella myndigheterna har fog för att i förekommande fall genomföra förhör för att bedöma fakta och omständigheter avseende den asylsökandes påstådda sexuella läggning, strider förhör om detaljer beträffande sökandens sexuella vanor mot de grundläggande rättigheter som säkerställs genom stadgan och framför allt mot rätten till respekt för privatlivet och familjelivet enligt artikel 7 i stadgan.
Vad därefter gäller möjligheten för de nationella myndigheterna att godta att, såsom har föreslagits av vissa av klagandena i de nationella målen, en asylsökande genomgår eventuella ”test” för fastställande av personens homosexuella läggning eller ger in bevis såsom videoupptagningar som visar när vederbörande utför intima handlingar, framhåller domstolen att förutom att sådan bevisning inte nödvändigtvis har något bevisvärde, kan den inkräkta på människans värdighet, som ska respekteras enligt artikel 1 i stadgan.
Att tillåta eller godta en sådan typ av bevisning skulle dessutom leda till en stimulanseffekt i förhållande till andra asylsökande och för dessa de facto innebära ett krav på att inge den typen av bevis.
När det gäller de behöriga myndigheternas möjlighet att göra bedömningen att den asylsökande brister i trovärdighet bland annat när sökanden inte åberopade sin påstådda sexuella läggning första gången han eller hon gavs tillfälle att lägga fram skälen till förföljelse, gör domstolen följande bedömning.
Det framgår av bestämmelserna i artikel 4.1 i direktiv 2004/83 att medlemsstaterna får betrakta det som den sökandes skyldighet att ”så snart som möjligt” lägga fram alla faktorer som behövs för att styrka ansökan om internationellt skydd.
Med hänsyn till att frågor som rör en persons personliga sfär, och framför allt en persons sexualitet, är känsliga till sin natur kan man dock inte dra slutsatsen att en person saknar trovärdighet endast därför att han eller hon på grund av sin tveksamhet att röja uppgifter om vissa intima aspekter av sitt liv inte omedelbart har berättat om sin homosexuella läggning.
Dessutom ska det påpekas att skyldigheten enligt artikel 4.1 i direktiv 2004/83 att ”så snart som möjligt” lägga fram alla faktorer som behövs för att styrka ansökan om internationellt skydd mildras av kravet på de behöriga myndigheterna enligt artikel 13.3 a direktiv 2005/85 och artikel 4.3 i direktiv 2004/83, att vid intervjun beakta de personliga och allmänna omständigheter som ligger bakom ansökan, inklusive sökandens utsatta ställning, och att göra en individuell bedömning av en ansökan samt beakta varje sökandes personliga ställning och förhållanden.
Att bedöma att en asylsökande brister i trovärdighet endast av det skälet att sökanden inte avslöjade sin sexuella läggning första gången han eller hon gavs tillfälle att lägga fram skälen till förföljelse skulle strida mot det i föregående punkt angivna kravet.
Mot bakgrund av det ovan anförda ska den fråga som har hänskjutits i vart och ett av målen C‑148/13–C‑150/13 bevaras enligt följande:
Artikel 4.3 c i direktiv 2004/83 samt artikel 13.3 a i direktiv 2005/85 ska tolkas så, att de utgör hinder för att de behöriga nationella myndigheterna, inom ramen för sin bedömning av fakta och omständigheter – som kan bli föremål för prövning i domstol – för att fastställa den sexuella läggningen hos en asylsökande, som till stöd för sin asylansökan har åberopat fruktan för förföljelse på grund av denna läggning, prövar den asylsökandes uppgifter och de skriftliga eller andra bevis som har åberopats till stöd för ansökan med hjälp av förhör som uteslutande baseras på stereotypa uppfattningar om homosexuella.
Artikel 4 i direktiv 2004/83, jämförd med artikel 7 i stadgan, ska tolkas så, att den utgör hinder för att de behöriga nationella myndigheterna, inom ramen för denna bedömning, genomför detaljerade förhör om den asylsökandes sexuella vanor.
Artikel 4 i direktiv 2004/83, jämförd med artikel 1 i stadgan, ska tolkas så, att den utgör hinder för att nämnda myndigheter, inom ramen för denna bedömning, såsom bevisning godtar att den asylsökande utför homosexuella handlingar, genomgår ”test” för fastställande av sin homosexuella läggning eller ger in videoupptagningar av homosexuella handlingar.
Artikel 4.3 i direktiv 2004/83 samt artikel 13.3 a i direktiv 2005/85 ska tolkas så, att de utgör hinder för att de behöriga nationella myndigheterna, inom ramen för samma bedömning, slår fast att den asylsökandes uppgifter brister i trovärdighet redan av det skälet att sökanden inte åberopade sin påstådda sexuella läggning första gången han eller hon gavs tillfälle att lägga fram skälen till förföljelse.
Rättegångskostnader
Eftersom förfarandet i förhållande till parterna i det nationella målet utgör ett led i beredningen av samma mål, ankommer det på den hänskjutande domstolen att besluta om rättegångskostnaderna. De kostnader för att avge yttrande till domstolen som andra än nämnda parter har haft är inte ersättningsgilla.
Mot denna bakgrund beslutar domstolen (stora avdelningen) följande:
Artikel 4.3 c i rådets direktiv 2004/83/EG av den 29 april 2004 om miniminormer för när tredjelandsmedborgare eller statslösa personer skall betraktas som flyktingar eller som personer som av andra skäl behöver internationellt skydd samt om dessa personers rättsliga ställning och om innehållet i det beviljade skyddet och artikel 13.3 a i rådets direktiv 2005/85/EG av den 1 december 2005 om miniminormer för medlemsstaternas förfaranden för beviljande eller återkallande av flyktingstatus ska tolkas så, att de utgör hinder för att de behöriga nationella myndigheterna, inom ramen för sin bedömning av fakta och omständigheter – som kan bli föremål för prövning i domstol – för att fastställa den sexuella läggningen hos en asylsökande, som till stöd för sin asylansökan har åberopat fruktan för förföljelse på grund av denna läggning, prövar den asylsökandes uppgifter och de skriftliga eller andra bevis som har åberopats till stöd för ansökan med hjälp av förhör som uteslutande baseras på stereotypa uppfattningar om homosexuella.
Artikel 4 i direktiv 2004/83, jämförd med artikel 7 i Europeiska unionens stadga om de grundläggande rättigheterna, ska tolkas så, att den utgör hinder för att de behöriga nationella myndigheterna, inom ramen för denna bedömning, genomför detaljerade förhör om den asylsökandes sexuella vanor.
Artikel 4 i direktiv 2004/83, jämförd med artikel 1 i Europeiska unionens stadga om de grundläggande rättigheterna, ska tolkas så, att den utgör hinder för att nämnda myndigheter, inom ramen för denna bedömning, såsom bevisning godtar att den asylsökande utför homosexuella handlingar, genomgår ”test” för fastställande av sin homosexuella läggning eller ger in videoupptagningar av homosexuella handlingar.
Artikel 4.3 i direktiv 2004/83 samt artikel 13.3 a i direktiv 2005/85 ska tolkas så, att de utgör hinder för att de behöriga nationella myndigheterna, inom ramen för samma bedömning, slår fast att den asylsökandes uppgifter brister i trovärdighet redan av det skälet att sökanden inte åberopade sin påstådda sexuella läggning första gången han eller hon gavs tillfälle att lägga fram skälen till förföljelse.
